module dct_comp (
    input wire clk,
    input wire rst_n,
    input wire [31:0] log_out,
    input wire log_valid,
    input wire [7:0] num_mfcc_coeffs,
    output reg [31:0] dct_out,
    output reg dct_valid
);

// Constants
localparam MAX_COEFFS = 32;

// DCT coefficients (stored in ROM)
reg [31:0] dct_coeffs [0:MAX_COEFFS-1][0:MAX_COEFFS-1];

// Intermediate variables
reg [31:0] dct_sum;
reg [$clog2(MAX_COEFFS)-1:0] coeff_idx;
reg [$clog2(MAX_COEFFS)-1:0] log_idx;

// DCT computation pipeline
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        dct_out <= 32'h0;
        dct_valid <= 1'b0;
        dct_sum <= 32'h0;
        coeff_idx <= 'h0;
        log_idx <= 'h0;
    end else if (log_valid) begin
        dct_sum <= dct_sum + (log_out * dct_coeffs[coeff_idx][log_idx]);
        log_idx <= log_idx + 1;

        if (log_idx == num_mfcc_coeffs - 1) begin
            dct_out <= dct_sum;
            dct_valid <= 1'b1;
            dct_sum <= 32'h0;
            coeff_idx <= coeff_idx + 1;
            log_idx <= 'h0;

            if (coeff_idx == num_mfcc_coeffs - 1) begin
                coeff_idx <= 'h0;
            end
        end else begin
            dct_valid <= 1'b0;
        end
    end else begin
        dct_valid <= 1'b0;
    end
end

// Initialize DCT coefficients 
initial begin
      dct_coeffs[0][0] = 32'h0B504F33;
      dct_coeffs[0][1] = 32'h0B504F33;
      dct_coeffs[0][2] = 32'h0B504F33;
      dct_coeffs[0][3] = 32'h0B504F33;
      dct_coeffs[0][4] = 32'h0B504F33;
      dct_coeffs[0][5] = 32'h0B504F33;
      dct_coeffs[0][6] = 32'h0B504F33;
      dct_coeffs[0][7] = 32'h0B504F33;
      dct_coeffs[0][8] = 32'h0B504F33;
      dct_coeffs[0][9] = 32'h0B504F33;
      dct_coeffs[0][10] = 32'h0B504F33;
      dct_coeffs[0][11] = 32'h0B504F33;
      dct_coeffs[0][12] = 32'h0B504F33;
      dct_coeffs[0][13] = 32'h0B504F33;
      dct_coeffs[0][14] = 32'h0B504F33;
      dct_coeffs[0][15] = 32'h0B504F33;
      dct_coeffs[0][16] = 32'h0B504F33;
      dct_coeffs[0][17] = 32'h0B504F33;
      dct_coeffs[0][18] = 32'h0B504F33;
      dct_coeffs[0][19] = 32'h0B504F33;
      dct_coeffs[0][20] = 32'h0B504F33;
      dct_coeffs[0][21] = 32'h0B504F33;
      dct_coeffs[0][22] = 32'h0B504F33;
      dct_coeffs[0][23] = 32'h0B504F33;
      dct_coeffs[0][24] = 32'h0B504F33;
      dct_coeffs[0][25] = 32'h0B504F33;
      dct_coeffs[0][26] = 32'h0B504F33;
      dct_coeffs[0][27] = 32'h0B504F33;
      dct_coeffs[0][28] = 32'h0B504F33;
      dct_coeffs[0][29] = 32'h0B504F33;
      dct_coeffs[0][30] = 32'h0B504F33;
      dct_coeffs[0][31] = 32'h0B504F33;
      dct_coeffs[1][0] = 32'h0FFB10F1;
      dct_coeffs[1][1] = 32'h0FD3AABF;
      dct_coeffs[1][2] = 32'h0F853F7D;
      dct_coeffs[1][3] = 32'h0F109082;
      dct_coeffs[1][4] = 32'h0E76BD7A;
      dct_coeffs[1][5] = 32'h0DB941A2;
      dct_coeffs[1][6] = 32'h0CD9F023;
      dct_coeffs[1][7] = 32'h0BDAEF91;
      dct_coeffs[1][8] = 32'h0ABEB49A;
      dct_coeffs[1][9] = 32'h0987FBFE;
      dct_coeffs[1][10] = 32'h0839C3CC;
      dct_coeffs[1][11] = 32'h06D74402;
      dct_coeffs[1][12] = 32'h0563E69D;
      dct_coeffs[1][13] = 32'h03E33F2F;
      dct_coeffs[1][14] = 32'h0259020D;
      dct_coeffs[1][15] = 32'h00C8FB2F;
      dct_coeffs[1][16] = 32'hFF3704D1;
      dct_coeffs[1][17] = 32'hFDA6FDF3;
      dct_coeffs[1][18] = 32'hFC1CC0D1;
      dct_coeffs[1][19] = 32'hFA9C1963;
      dct_coeffs[1][20] = 32'hF928BBFE;
      dct_coeffs[1][21] = 32'hF7C63C34;
      dct_coeffs[1][22] = 32'hF6780402;
      dct_coeffs[1][23] = 32'hF5414B66;
      dct_coeffs[1][24] = 32'hF425106F;
      dct_coeffs[1][25] = 32'hF3260FDD;
      dct_coeffs[1][26] = 32'hF246BE5E;
      dct_coeffs[1][27] = 32'hF1894286;
      dct_coeffs[1][28] = 32'hF0EF6F7E;
      dct_coeffs[1][29] = 32'hF07AC083;
      dct_coeffs[1][30] = 32'hF02C5541;
      dct_coeffs[1][31] = 32'hF004EF0F;
      dct_coeffs[2][0] = 32'h0FEC46D1;
      dct_coeffs[2][1] = 32'h0F4FA0AB;
      dct_coeffs[2][2] = 32'h0E1C5978;
      dct_coeffs[2][3] = 32'h0C5E4035;
      dct_coeffs[2][4] = 32'h0A267992;
      dct_coeffs[2][5] = 32'h078AD74E;
      dct_coeffs[2][6] = 32'h04A5018B;
      dct_coeffs[2][7] = 32'h01917A6B;
      dct_coeffs[2][8] = 32'hFE6E8595;
      dct_coeffs[2][9] = 32'hFB5AFE75;
      dct_coeffs[2][10] = 32'hF87528B2;
      dct_coeffs[2][11] = 32'hF5D9866E;
      dct_coeffs[2][12] = 32'hF3A1BFCB;
      dct_coeffs[2][13] = 32'hF1E3A688;
      dct_coeffs[2][14] = 32'hF0B05F55;
      dct_coeffs[2][15] = 32'hF013B92F;
      dct_coeffs[2][16] = 32'hF013B92F;
      dct_coeffs[2][17] = 32'hF0B05F55;
      dct_coeffs[2][18] = 32'hF1E3A688;
      dct_coeffs[2][19] = 32'hF3A1BFCB;
      dct_coeffs[2][20] = 32'hF5D9866E;
      dct_coeffs[2][21] = 32'hF87528B2;
      dct_coeffs[2][22] = 32'hFB5AFE75;
      dct_coeffs[2][23] = 32'hFE6E8595;
      dct_coeffs[2][24] = 32'h01917A6B;
      dct_coeffs[2][25] = 32'h04A5018B;
      dct_coeffs[2][26] = 32'h078AD74E;
      dct_coeffs[2][27] = 32'h0A267992;
      dct_coeffs[2][28] = 32'h0C5E4035;
      dct_coeffs[2][29] = 32'h0E1C5978;
      dct_coeffs[2][30] = 32'h0F4FA0AB;
      dct_coeffs[2][31] = 32'h0FEC46D1;
      dct_coeffs[3][0] = 32'h0FD3AABF;
      dct_coeffs[3][1] = 32'h0E76BD7A;
      dct_coeffs[3][2] = 32'h0BDAEF91;
      dct_coeffs[3][3] = 32'h0839C3CC;
      dct_coeffs[3][4] = 32'h03E33F2F;
      dct_coeffs[3][5] = 32'hFF3704D1;
      dct_coeffs[3][6] = 32'hFA9C1963;
      dct_coeffs[3][7] = 32'hF6780402;
      dct_coeffs[3][8] = 32'hF3260FDD;
      dct_coeffs[3][9] = 32'hF0EF6F7E;
      dct_coeffs[3][10] = 32'hF004EF0F;
      dct_coeffs[3][11] = 32'hF07AC083;
      dct_coeffs[3][12] = 32'hF246BE5E;
      dct_coeffs[3][13] = 32'hF5414B66;
      dct_coeffs[3][14] = 32'hF928BBFE;
      dct_coeffs[3][15] = 32'hFDA6FDF3;
      dct_coeffs[3][16] = 32'h0259020D;
      dct_coeffs[3][17] = 32'h06D74402;
      dct_coeffs[3][18] = 32'h0ABEB49A;
      dct_coeffs[3][19] = 32'h0DB941A2;
      dct_coeffs[3][20] = 32'h0F853F7D;
      dct_coeffs[3][21] = 32'h0FFB10F1;
      dct_coeffs[3][22] = 32'h0F109082;
      dct_coeffs[3][23] = 32'h0CD9F023;
      dct_coeffs[3][24] = 32'h0987FBFE;
      dct_coeffs[3][25] = 32'h0563E69D;
      dct_coeffs[3][26] = 32'h00C8FB2F;
      dct_coeffs[3][27] = 32'hFC1CC0D1;
      dct_coeffs[3][28] = 32'hF7C63C34;
      dct_coeffs[3][29] = 32'hF425106F;
      dct_coeffs[3][30] = 32'hF1894286;
      dct_coeffs[3][31] = 32'hF02C5541;
      dct_coeffs[4][0] = 32'h0FB14BE7;
      dct_coeffs[4][1] = 32'h0D4DB314;
      dct_coeffs[4][2] = 32'h08E39D9C;
      dct_coeffs[4][3] = 32'h031F1707;
      dct_coeffs[4][4] = 32'hFCE0E8F9;
      dct_coeffs[4][5] = 32'hF71C6264;
      dct_coeffs[4][6] = 32'hF2B24CEC;
      dct_coeffs[4][7] = 32'hF04EB419;
      dct_coeffs[4][8] = 32'hF04EB419;
      dct_coeffs[4][9] = 32'hF2B24CEC;
      dct_coeffs[4][10] = 32'hF71C6264;
      dct_coeffs[4][11] = 32'hFCE0E8F9;
      dct_coeffs[4][12] = 32'h031F1707;
      dct_coeffs[4][13] = 32'h08E39D9C;
      dct_coeffs[4][14] = 32'h0D4DB314;
      dct_coeffs[4][15] = 32'h0FB14BE7;
      dct_coeffs[4][16] = 32'h0FB14BE7;
      dct_coeffs[4][17] = 32'h0D4DB314;
      dct_coeffs[4][18] = 32'h08E39D9C;
      dct_coeffs[4][19] = 32'h031F1707;
      dct_coeffs[4][20] = 32'hFCE0E8F9;
      dct_coeffs[4][21] = 32'hF71C6264;
      dct_coeffs[4][22] = 32'hF2B24CEC;
      dct_coeffs[4][23] = 32'hF04EB419;
      dct_coeffs[4][24] = 32'hF04EB419;
      dct_coeffs[4][25] = 32'hF2B24CEC;
      dct_coeffs[4][26] = 32'hF71C6264;
      dct_coeffs[4][27] = 32'hFCE0E8F9;
      dct_coeffs[4][28] = 32'h031F1707;
      dct_coeffs[4][29] = 32'h08E39D9C;
      dct_coeffs[4][30] = 32'h0D4DB314;
      dct_coeffs[4][31] = 32'h0FB14BE7;
      dct_coeffs[5][0] = 32'h0F853F7D;
      dct_coeffs[5][1] = 32'h0BDAEF91;
      dct_coeffs[5][2] = 32'h0563E69D;
      dct_coeffs[5][3] = 32'hFDA6FDF3;
      dct_coeffs[5][4] = 32'hF6780402;
      dct_coeffs[5][5] = 32'hF1894286;
      dct_coeffs[5][6] = 32'hF004EF0F;
      dct_coeffs[5][7] = 32'hF246BE5E;
      dct_coeffs[5][8] = 32'hF7C63C34;
      dct_coeffs[5][9] = 32'hFF3704D1;
      dct_coeffs[5][10] = 32'h06D74402;
      dct_coeffs[5][11] = 32'h0CD9F023;
      dct_coeffs[5][12] = 32'h0FD3AABF;
      dct_coeffs[5][13] = 32'h0F109082;
      dct_coeffs[5][14] = 32'h0ABEB49A;
      dct_coeffs[5][15] = 32'h03E33F2F;
      dct_coeffs[5][16] = 32'hFC1CC0D1;
      dct_coeffs[5][17] = 32'hF5414B66;
      dct_coeffs[5][18] = 32'hF0EF6F7E;
      dct_coeffs[5][19] = 32'hF02C5541;
      dct_coeffs[5][20] = 32'hF3260FDD;
      dct_coeffs[5][21] = 32'hF928BBFE;
      dct_coeffs[5][22] = 32'h00C8FB2F;
      dct_coeffs[5][23] = 32'h0839C3CC;
      dct_coeffs[5][24] = 32'h0DB941A2;
      dct_coeffs[5][25] = 32'h0FFB10F1;
      dct_coeffs[5][26] = 32'h0E76BD7A;
      dct_coeffs[5][27] = 32'h0987FBFE;
      dct_coeffs[5][28] = 32'h0259020D;
      dct_coeffs[5][29] = 32'hFA9C1963;
      dct_coeffs[5][30] = 32'hF425106F;
      dct_coeffs[5][31] = 32'hF07AC083;
      dct_coeffs[6][0] = 32'h0F4FA0AB;
      dct_coeffs[6][1] = 32'h0A267992;
      dct_coeffs[6][2] = 32'h01917A6B;
      dct_coeffs[6][3] = 32'hF87528B2;
      dct_coeffs[6][4] = 32'hF1E3A688;
      dct_coeffs[6][5] = 32'hF013B92F;
      dct_coeffs[6][6] = 32'hF3A1BFCB;
      dct_coeffs[6][7] = 32'hFB5AFE75;
      dct_coeffs[6][8] = 32'h04A5018B;
      dct_coeffs[6][9] = 32'h0C5E4035;
      dct_coeffs[6][10] = 32'h0FEC46D1;
      dct_coeffs[6][11] = 32'h0E1C5978;
      dct_coeffs[6][12] = 32'h078AD74E;
      dct_coeffs[6][13] = 32'hFE6E8595;
      dct_coeffs[6][14] = 32'hF5D9866E;
      dct_coeffs[6][15] = 32'hF0B05F55;
      dct_coeffs[6][16] = 32'hF0B05F55;
      dct_coeffs[6][17] = 32'hF5D9866E;
      dct_coeffs[6][18] = 32'hFE6E8595;
      dct_coeffs[6][19] = 32'h078AD74E;
      dct_coeffs[6][20] = 32'h0E1C5978;
      dct_coeffs[6][21] = 32'h0FEC46D1;
      dct_coeffs[6][22] = 32'h0C5E4035;
      dct_coeffs[6][23] = 32'h04A5018B;
      dct_coeffs[6][24] = 32'hFB5AFE75;
      dct_coeffs[6][25] = 32'hF3A1BFCB;
      dct_coeffs[6][26] = 32'hF013B92F;
      dct_coeffs[6][27] = 32'hF1E3A688;
      dct_coeffs[6][28] = 32'hF87528B2;
      dct_coeffs[6][29] = 32'h01917A6B;
      dct_coeffs[6][30] = 32'h0A267992;
      dct_coeffs[6][31] = 32'h0F4FA0AB;
      dct_coeffs[7][0] = 32'h0F109082;
      dct_coeffs[7][1] = 32'h0839C3CC;
      dct_coeffs[7][2] = 32'hFDA6FDF3;
      dct_coeffs[7][3] = 32'hF425106F;
      dct_coeffs[7][4] = 32'hF004EF0F;
      dct_coeffs[7][5] = 32'hF3260FDD;
      dct_coeffs[7][6] = 32'hFC1CC0D1;
      dct_coeffs[7][7] = 32'h06D74402;
      dct_coeffs[7][8] = 32'h0E76BD7A;
      dct_coeffs[7][9] = 32'h0F853F7D;
      dct_coeffs[7][10] = 32'h0987FBFE;
      dct_coeffs[7][11] = 32'hFF3704D1;
      dct_coeffs[7][12] = 32'hF5414B66;
      dct_coeffs[7][13] = 32'hF02C5541;
      dct_coeffs[7][14] = 32'hF246BE5E;
      dct_coeffs[7][15] = 32'hFA9C1963;
      dct_coeffs[7][16] = 32'h0563E69D;
      dct_coeffs[7][17] = 32'h0DB941A2;
      dct_coeffs[7][18] = 32'h0FD3AABF;
      dct_coeffs[7][19] = 32'h0ABEB49A;
      dct_coeffs[7][20] = 32'h00C8FB2F;
      dct_coeffs[7][21] = 32'hF6780402;
      dct_coeffs[7][22] = 32'hF07AC083;
      dct_coeffs[7][23] = 32'hF1894286;
      dct_coeffs[7][24] = 32'hF928BBFE;
      dct_coeffs[7][25] = 32'h03E33F2F;
      dct_coeffs[7][26] = 32'h0CD9F023;
      dct_coeffs[7][27] = 32'h0FFB10F1;
      dct_coeffs[7][28] = 32'h0BDAEF91;
      dct_coeffs[7][29] = 32'h0259020D;
      dct_coeffs[7][30] = 32'hF7C63C34;
      dct_coeffs[7][31] = 32'hF0EF6F7E;
      dct_coeffs[8][0] = 32'h0EC835E7;
      dct_coeffs[8][1] = 32'h061F78A9;
      dct_coeffs[8][2] = 32'hF9E08757;
      dct_coeffs[8][3] = 32'hF137CA19;
      dct_coeffs[8][4] = 32'hF137CA19;
      dct_coeffs[8][5] = 32'hF9E08757;
      dct_coeffs[8][6] = 32'h061F78A9;
      dct_coeffs[8][7] = 32'h0EC835E7;
      dct_coeffs[8][8] = 32'h0EC835E7;
      dct_coeffs[8][9] = 32'h061F78A9;
      dct_coeffs[8][10] = 32'hF9E08757;
      dct_coeffs[8][11] = 32'hF137CA19;
      dct_coeffs[8][12] = 32'hF137CA19;
      dct_coeffs[8][13] = 32'hF9E08757;
      dct_coeffs[8][14] = 32'h061F78A9;
      dct_coeffs[8][15] = 32'h0EC835E7;
      dct_coeffs[8][16] = 32'h0EC835E7;
      dct_coeffs[8][17] = 32'h061F78A9;
      dct_coeffs[8][18] = 32'hF9E08757;
      dct_coeffs[8][19] = 32'hF137CA19;
      dct_coeffs[8][20] = 32'hF137CA19;
      dct_coeffs[8][21] = 32'hF9E08757;
      dct_coeffs[8][22] = 32'h061F78A9;
      dct_coeffs[8][23] = 32'h0EC835E7;
      dct_coeffs[8][24] = 32'h0EC835E7;
      dct_coeffs[8][25] = 32'h061F78A9;
      dct_coeffs[8][26] = 32'hF9E08757;
      dct_coeffs[8][27] = 32'hF137CA19;
      dct_coeffs[8][28] = 32'hF137CA19;
      dct_coeffs[8][29] = 32'hF9E08757;
      dct_coeffs[8][30] = 32'h061F78A9;
      dct_coeffs[8][31] = 32'h0EC835E7;
      dct_coeffs[9][0] = 32'h0E76BD7A;
      dct_coeffs[9][1] = 32'h03E33F2F;
      dct_coeffs[9][2] = 32'hF6780402;
      dct_coeffs[9][3] = 32'hF004EF0F;
      dct_coeffs[9][4] = 32'hF5414B66;
      dct_coeffs[9][5] = 32'h0259020D;
      dct_coeffs[9][6] = 32'h0DB941A2;
      dct_coeffs[9][7] = 32'h0F109082;
      dct_coeffs[9][8] = 32'h0563E69D;
      dct_coeffs[9][9] = 32'hF7C63C34;
      dct_coeffs[9][10] = 32'hF02C5541;
      dct_coeffs[9][11] = 32'hF425106F;
      dct_coeffs[9][12] = 32'h00C8FB2F;
      dct_coeffs[9][13] = 32'h0CD9F023;
      dct_coeffs[9][14] = 32'h0F853F7D;
      dct_coeffs[9][15] = 32'h06D74402;
      dct_coeffs[9][16] = 32'hF928BBFE;
      dct_coeffs[9][17] = 32'hF07AC083;
      dct_coeffs[9][18] = 32'hF3260FDD;
      dct_coeffs[9][19] = 32'hFF3704D1;
      dct_coeffs[9][20] = 32'h0BDAEF91;
      dct_coeffs[9][21] = 32'h0FD3AABF;
      dct_coeffs[9][22] = 32'h0839C3CC;
      dct_coeffs[9][23] = 32'hFA9C1963;
      dct_coeffs[9][24] = 32'hF0EF6F7E;
      dct_coeffs[9][25] = 32'hF246BE5E;
      dct_coeffs[9][26] = 32'hFDA6FDF3;
      dct_coeffs[9][27] = 32'h0ABEB49A;
      dct_coeffs[9][28] = 32'h0FFB10F1;
      dct_coeffs[9][29] = 32'h0987FBFE;
      dct_coeffs[9][30] = 32'hFC1CC0D1;
      dct_coeffs[9][31] = 32'hF1894286;
      dct_coeffs[10][0] = 32'h0E1C5978;
      dct_coeffs[10][1] = 32'h01917A6B;
      dct_coeffs[10][2] = 32'hF3A1BFCB;
      dct_coeffs[10][3] = 32'hF0B05F55;
      dct_coeffs[10][4] = 32'hFB5AFE75;
      dct_coeffs[10][5] = 32'h0A267992;
      dct_coeffs[10][6] = 32'h0FEC46D1;
      dct_coeffs[10][7] = 32'h078AD74E;
      dct_coeffs[10][8] = 32'hF87528B2;
      dct_coeffs[10][9] = 32'hF013B92F;
      dct_coeffs[10][10] = 32'hF5D9866E;
      dct_coeffs[10][11] = 32'h04A5018B;
      dct_coeffs[10][12] = 32'h0F4FA0AB;
      dct_coeffs[10][13] = 32'h0C5E4035;
      dct_coeffs[10][14] = 32'hFE6E8595;
      dct_coeffs[10][15] = 32'hF1E3A688;
      dct_coeffs[10][16] = 32'hF1E3A688;
      dct_coeffs[10][17] = 32'hFE6E8595;
      dct_coeffs[10][18] = 32'h0C5E4035;
      dct_coeffs[10][19] = 32'h0F4FA0AB;
      dct_coeffs[10][20] = 32'h04A5018B;
      dct_coeffs[10][21] = 32'hF5D9866E;
      dct_coeffs[10][22] = 32'hF013B92F;
      dct_coeffs[10][23] = 32'hF87528B2;
      dct_coeffs[10][24] = 32'h078AD74E;
      dct_coeffs[10][25] = 32'h0FEC46D1;
      dct_coeffs[10][26] = 32'h0A267992;
      dct_coeffs[10][27] = 32'hFB5AFE75;
      dct_coeffs[10][28] = 32'hF0B05F55;
      dct_coeffs[10][29] = 32'hF3A1BFCB;
      dct_coeffs[10][30] = 32'h01917A6B;
      dct_coeffs[10][31] = 32'h0E1C5978;
      dct_coeffs[11][0] = 32'h0DB941A2;
      dct_coeffs[11][1] = 32'hFF3704D1;
      dct_coeffs[11][2] = 32'hF1894286;
      dct_coeffs[11][3] = 32'hF3260FDD;
      dct_coeffs[11][4] = 32'h0259020D;
      dct_coeffs[11][5] = 32'h0F109082;
      dct_coeffs[11][6] = 32'h0BDAEF91;
      dct_coeffs[11][7] = 32'hFC1CC0D1;
      dct_coeffs[11][8] = 32'hF07AC083;
      dct_coeffs[11][9] = 32'hF5414B66;
      dct_coeffs[11][10] = 32'h0563E69D;
      dct_coeffs[11][11] = 32'h0FD3AABF;
      dct_coeffs[11][12] = 32'h0987FBFE;
      dct_coeffs[11][13] = 32'hF928BBFE;
      dct_coeffs[11][14] = 32'hF004EF0F;
      dct_coeffs[11][15] = 32'hF7C63C34;
      dct_coeffs[11][16] = 32'h0839C3CC;
      dct_coeffs[11][17] = 32'h0FFB10F1;
      dct_coeffs[11][18] = 32'h06D74402;
      dct_coeffs[11][19] = 32'hF6780402;
      dct_coeffs[11][20] = 32'hF02C5541;
      dct_coeffs[11][21] = 32'hFA9C1963;
      dct_coeffs[11][22] = 32'h0ABEB49A;
      dct_coeffs[11][23] = 32'h0F853F7D;
      dct_coeffs[11][24] = 32'h03E33F2F;
      dct_coeffs[11][25] = 32'hF425106F;
      dct_coeffs[11][26] = 32'hF0EF6F7E;
      dct_coeffs[11][27] = 32'hFDA6FDF3;
      dct_coeffs[11][28] = 32'h0CD9F023;
      dct_coeffs[11][29] = 32'h0E76BD7A;
      dct_coeffs[11][30] = 32'h00C8FB2F;
      dct_coeffs[11][31] = 32'hF246BE5E;
      dct_coeffs[12][0] = 32'h0D4DB314;
      dct_coeffs[12][1] = 32'hFCE0E8F9;
      dct_coeffs[12][2] = 32'hF04EB419;
      dct_coeffs[12][3] = 32'hF71C6264;
      dct_coeffs[12][4] = 32'h08E39D9C;
      dct_coeffs[12][5] = 32'h0FB14BE7;
      dct_coeffs[12][6] = 32'h031F1707;
      dct_coeffs[12][7] = 32'hF2B24CEC;
      dct_coeffs[12][8] = 32'hF2B24CEC;
      dct_coeffs[12][9] = 32'h031F1707;
      dct_coeffs[12][10] = 32'h0FB14BE7;
      dct_coeffs[12][11] = 32'h08E39D9C;
      dct_coeffs[12][12] = 32'hF71C6264;
      dct_coeffs[12][13] = 32'hF04EB419;
      dct_coeffs[12][14] = 32'hFCE0E8F9;
      dct_coeffs[12][15] = 32'h0D4DB314;
      dct_coeffs[12][16] = 32'h0D4DB314;
      dct_coeffs[12][17] = 32'hFCE0E8F9;
      dct_coeffs[12][18] = 32'hF04EB419;
      dct_coeffs[12][19] = 32'hF71C6264;
      dct_coeffs[12][20] = 32'h08E39D9C;
      dct_coeffs[12][21] = 32'h0FB14BE7;
      dct_coeffs[12][22] = 32'h031F1707;
      dct_coeffs[12][23] = 32'hF2B24CEC;
      dct_coeffs[12][24] = 32'hF2B24CEC;
      dct_coeffs[12][25] = 32'h031F1707;
      dct_coeffs[12][26] = 32'h0FB14BE7;
      dct_coeffs[12][27] = 32'h08E39D9C;
      dct_coeffs[12][28] = 32'hF71C6264;
      dct_coeffs[12][29] = 32'hF04EB419;
      dct_coeffs[12][30] = 32'hFCE0E8F9;
      dct_coeffs[12][31] = 32'h0D4DB314;
      dct_coeffs[13][0] = 32'h0CD9F023;
      dct_coeffs[13][1] = 32'hFA9C1963;
      dct_coeffs[13][2] = 32'hF004EF0F;
      dct_coeffs[13][3] = 32'hFC1CC0D1;
      dct_coeffs[13][4] = 32'h0DB941A2;
      dct_coeffs[13][5] = 32'h0BDAEF91;
      dct_coeffs[13][6] = 32'hF928BBFE;
      dct_coeffs[13][7] = 32'hF02C5541;
      dct_coeffs[13][8] = 32'hFDA6FDF3;
      dct_coeffs[13][9] = 32'h0E76BD7A;
      dct_coeffs[13][10] = 32'h0ABEB49A;
      dct_coeffs[13][11] = 32'hF7C63C34;
      dct_coeffs[13][12] = 32'hF07AC083;
      dct_coeffs[13][13] = 32'hFF3704D1;
      dct_coeffs[13][14] = 32'h0F109082;
      dct_coeffs[13][15] = 32'h0987FBFE;
      dct_coeffs[13][16] = 32'hF6780402;
      dct_coeffs[13][17] = 32'hF0EF6F7E;
      dct_coeffs[13][18] = 32'h00C8FB2F;
      dct_coeffs[13][19] = 32'h0F853F7D;
      dct_coeffs[13][20] = 32'h0839C3CC;
      dct_coeffs[13][21] = 32'hF5414B66;
      dct_coeffs[13][22] = 32'hF1894286;
      dct_coeffs[13][23] = 32'h0259020D;
      dct_coeffs[13][24] = 32'h0FD3AABF;
      dct_coeffs[13][25] = 32'h06D74402;
      dct_coeffs[13][26] = 32'hF425106F;
      dct_coeffs[13][27] = 32'hF246BE5E;
      dct_coeffs[13][28] = 32'h03E33F2F;
      dct_coeffs[13][29] = 32'h0FFB10F1;
      dct_coeffs[13][30] = 32'h0563E69D;
      dct_coeffs[13][31] = 32'hF3260FDD;
      dct_coeffs[14][0] = 32'h0C5E4035;
      dct_coeffs[14][1] = 32'hF87528B2;
      dct_coeffs[14][2] = 32'hF0B05F55;
      dct_coeffs[14][3] = 32'h01917A6B;
      dct_coeffs[14][4] = 32'h0FEC46D1;
      dct_coeffs[14][5] = 32'h04A5018B;
      dct_coeffs[14][6] = 32'hF1E3A688;
      dct_coeffs[14][7] = 32'hF5D9866E;
      dct_coeffs[14][8] = 32'h0A267992;
      dct_coeffs[14][9] = 32'h0E1C5978;
      dct_coeffs[14][10] = 32'hFB5AFE75;
      dct_coeffs[14][11] = 32'hF013B92F;
      dct_coeffs[14][12] = 32'hFE6E8595;
      dct_coeffs[14][13] = 32'h0F4FA0AB;
      dct_coeffs[14][14] = 32'h078AD74E;
      dct_coeffs[14][15] = 32'hF3A1BFCB;
      dct_coeffs[14][16] = 32'hF3A1BFCB;
      dct_coeffs[14][17] = 32'h078AD74E;
      dct_coeffs[14][18] = 32'h0F4FA0AB;
      dct_coeffs[14][19] = 32'hFE6E8595;
      dct_coeffs[14][20] = 32'hF013B92F;
      dct_coeffs[14][21] = 32'hFB5AFE75;
      dct_coeffs[14][22] = 32'h0E1C5978;
      dct_coeffs[14][23] = 32'h0A267992;
      dct_coeffs[14][24] = 32'hF5D9866E;
      dct_coeffs[14][25] = 32'hF1E3A688;
      dct_coeffs[14][26] = 32'h04A5018B;
      dct_coeffs[14][27] = 32'h0FEC46D1;
      dct_coeffs[14][28] = 32'h01917A6B;
      dct_coeffs[14][29] = 32'hF0B05F55;
      dct_coeffs[14][30] = 32'hF87528B2;
      dct_coeffs[14][31] = 32'h0C5E4035;
      dct_coeffs[15][0] = 32'h0BDAEF91;
      dct_coeffs[15][1] = 32'hF6780402;
      dct_coeffs[15][2] = 32'hF246BE5E;
      dct_coeffs[15][3] = 32'h06D74402;
      dct_coeffs[15][4] = 32'h0F109082;
      dct_coeffs[15][5] = 32'hFC1CC0D1;
      dct_coeffs[15][6] = 32'hF02C5541;
      dct_coeffs[15][7] = 32'h00C8FB2F;
      dct_coeffs[15][8] = 32'h0FFB10F1;
      dct_coeffs[15][9] = 32'h0259020D;
      dct_coeffs[15][10] = 32'hF07AC083;
      dct_coeffs[15][11] = 32'hFA9C1963;
      dct_coeffs[15][12] = 32'h0E76BD7A;
      dct_coeffs[15][13] = 32'h0839C3CC;
      dct_coeffs[15][14] = 32'hF3260FDD;
      dct_coeffs[15][15] = 32'hF5414B66;
      dct_coeffs[15][16] = 32'h0ABEB49A;
      dct_coeffs[15][17] = 32'h0CD9F023;
      dct_coeffs[15][18] = 32'hF7C63C34;
      dct_coeffs[15][19] = 32'hF1894286;
      dct_coeffs[15][20] = 32'h0563E69D;
      dct_coeffs[15][21] = 32'h0F853F7D;
      dct_coeffs[15][22] = 32'hFDA6FDF3;
      dct_coeffs[15][23] = 32'hF004EF0F;
      dct_coeffs[15][24] = 32'hFF3704D1;
      dct_coeffs[15][25] = 32'h0FD3AABF;
      dct_coeffs[15][26] = 32'h03E33F2F;
      dct_coeffs[15][27] = 32'hF0EF6F7E;
      dct_coeffs[15][28] = 32'hF928BBFE;
      dct_coeffs[15][29] = 32'h0DB941A2;
      dct_coeffs[15][30] = 32'h0987FBFE;
      dct_coeffs[15][31] = 32'hF425106F;
      dct_coeffs[16][0] = 32'h0B504F33;
      dct_coeffs[16][1] = 32'hF4AFB0CD;
      dct_coeffs[16][2] = 32'hF4AFB0CD;
      dct_coeffs[16][3] = 32'h0B504F33;
      dct_coeffs[16][4] = 32'h0B504F33;
      dct_coeffs[16][5] = 32'hF4AFB0CD;
      dct_coeffs[16][6] = 32'hF4AFB0CD;
      dct_coeffs[16][7] = 32'h0B504F33;
      dct_coeffs[16][8] = 32'h0B504F33;
      dct_coeffs[16][9] = 32'hF4AFB0CD;
      dct_coeffs[16][10] = 32'hF4AFB0CD;
      dct_coeffs[16][11] = 32'h0B504F33;
      dct_coeffs[16][12] = 32'h0B504F33;
      dct_coeffs[16][13] = 32'hF4AFB0CD;
      dct_coeffs[16][14] = 32'hF4AFB0CD;
      dct_coeffs[16][15] = 32'h0B504F33;
      dct_coeffs[16][16] = 32'h0B504F33;
      dct_coeffs[16][17] = 32'hF4AFB0CD;
      dct_coeffs[16][18] = 32'hF4AFB0CD;
      dct_coeffs[16][19] = 32'h0B504F33;
      dct_coeffs[16][20] = 32'h0B504F33;
      dct_coeffs[16][21] = 32'hF4AFB0CD;
      dct_coeffs[16][22] = 32'hF4AFB0CD;
      dct_coeffs[16][23] = 32'h0B504F33;
      dct_coeffs[16][24] = 32'h0B504F33;
      dct_coeffs[16][25] = 32'hF4AFB0CD;
      dct_coeffs[16][26] = 32'hF4AFB0CD;
      dct_coeffs[16][27] = 32'h0B504F33;
      dct_coeffs[16][28] = 32'h0B504F33;
      dct_coeffs[16][29] = 32'hF4AFB0CD;
      dct_coeffs[16][30] = 32'hF4AFB0CD;
      dct_coeffs[16][31] = 32'h0B504F33;
      dct_coeffs[17][0] = 32'h0ABEB49A;
      dct_coeffs[17][1] = 32'hF3260FDD;
      dct_coeffs[17][2] = 32'hF7C63C34;
      dct_coeffs[17][3] = 32'h0E76BD7A;
      dct_coeffs[17][4] = 32'h0563E69D;
      dct_coeffs[17][5] = 32'hF07AC083;
      dct_coeffs[17][6] = 32'hFDA6FDF3;
      dct_coeffs[17][7] = 32'h0FFB10F1;
      dct_coeffs[17][8] = 32'hFF3704D1;
      dct_coeffs[17][9] = 32'hF02C5541;
      dct_coeffs[17][10] = 32'h03E33F2F;
      dct_coeffs[17][11] = 32'h0F109082;
      dct_coeffs[17][12] = 32'hF928BBFE;
      dct_coeffs[17][13] = 32'hF246BE5E;
      dct_coeffs[17][14] = 32'h0987FBFE;
      dct_coeffs[17][15] = 32'h0BDAEF91;
      dct_coeffs[17][16] = 32'hF425106F;
      dct_coeffs[17][17] = 32'hF6780402;
      dct_coeffs[17][18] = 32'h0DB941A2;
      dct_coeffs[17][19] = 32'h06D74402;
      dct_coeffs[17][20] = 32'hF0EF6F7E;
      dct_coeffs[17][21] = 32'hFC1CC0D1;
      dct_coeffs[17][22] = 32'h0FD3AABF;
      dct_coeffs[17][23] = 32'h00C8FB2F;
      dct_coeffs[17][24] = 32'hF004EF0F;
      dct_coeffs[17][25] = 32'h0259020D;
      dct_coeffs[17][26] = 32'h0F853F7D;
      dct_coeffs[17][27] = 32'hFA9C1963;
      dct_coeffs[17][28] = 32'hF1894286;
      dct_coeffs[17][29] = 32'h0839C3CC;
      dct_coeffs[17][30] = 32'h0CD9F023;
      dct_coeffs[17][31] = 32'hF5414B66;
      dct_coeffs[18][0] = 32'h0A267992;
      dct_coeffs[18][1] = 32'hF1E3A688;
      dct_coeffs[18][2] = 32'hFB5AFE75;
      dct_coeffs[18][3] = 32'h0FEC46D1;
      dct_coeffs[18][4] = 32'hFE6E8595;
      dct_coeffs[18][5] = 32'hF0B05F55;
      dct_coeffs[18][6] = 32'h078AD74E;
      dct_coeffs[18][7] = 32'h0C5E4035;
      dct_coeffs[18][8] = 32'hF3A1BFCB;
      dct_coeffs[18][9] = 32'hF87528B2;
      dct_coeffs[18][10] = 32'h0F4FA0AB;
      dct_coeffs[18][11] = 32'h01917A6B;
      dct_coeffs[18][12] = 32'hF013B92F;
      dct_coeffs[18][13] = 32'h04A5018B;
      dct_coeffs[18][14] = 32'h0E1C5978;
      dct_coeffs[18][15] = 32'hF5D9866E;
      dct_coeffs[18][16] = 32'hF5D9866E;
      dct_coeffs[18][17] = 32'h0E1C5978;
      dct_coeffs[18][18] = 32'h04A5018B;
      dct_coeffs[18][19] = 32'hF013B92F;
      dct_coeffs[18][20] = 32'h01917A6B;
      dct_coeffs[18][21] = 32'h0F4FA0AB;
      dct_coeffs[18][22] = 32'hF87528B2;
      dct_coeffs[18][23] = 32'hF3A1BFCB;
      dct_coeffs[18][24] = 32'h0C5E4035;
      dct_coeffs[18][25] = 32'h078AD74E;
      dct_coeffs[18][26] = 32'hF0B05F55;
      dct_coeffs[18][27] = 32'hFE6E8595;
      dct_coeffs[18][28] = 32'h0FEC46D1;
      dct_coeffs[18][29] = 32'hFB5AFE75;
      dct_coeffs[18][30] = 32'hF1E3A688;
      dct_coeffs[18][31] = 32'h0A267992;
      dct_coeffs[19][0] = 32'h0987FBFE;
      dct_coeffs[19][1] = 32'hF0EF6F7E;
      dct_coeffs[19][2] = 32'hFF3704D1;
      dct_coeffs[19][3] = 32'h0F853F7D;
      dct_coeffs[19][4] = 32'hF7C63C34;
      dct_coeffs[19][5] = 32'hF5414B66;
      dct_coeffs[19][6] = 32'h0E76BD7A;
      dct_coeffs[19][7] = 32'h0259020D;
      dct_coeffs[19][8] = 32'hF02C5541;
      dct_coeffs[19][9] = 32'h06D74402;
      dct_coeffs[19][10] = 32'h0BDAEF91;
      dct_coeffs[19][11] = 32'hF246BE5E;
      dct_coeffs[19][12] = 32'hFC1CC0D1;
      dct_coeffs[19][13] = 32'h0FFB10F1;
      dct_coeffs[19][14] = 32'hFA9C1963;
      dct_coeffs[19][15] = 32'hF3260FDD;
      dct_coeffs[19][16] = 32'h0CD9F023;
      dct_coeffs[19][17] = 32'h0563E69D;
      dct_coeffs[19][18] = 32'hF004EF0F;
      dct_coeffs[19][19] = 32'h03E33F2F;
      dct_coeffs[19][20] = 32'h0DB941A2;
      dct_coeffs[19][21] = 32'hF425106F;
      dct_coeffs[19][22] = 32'hF928BBFE;
      dct_coeffs[19][23] = 32'h0FD3AABF;
      dct_coeffs[19][24] = 32'hFDA6FDF3;
      dct_coeffs[19][25] = 32'hF1894286;
      dct_coeffs[19][26] = 32'h0ABEB49A;
      dct_coeffs[19][27] = 32'h0839C3CC;
      dct_coeffs[19][28] = 32'hF07AC083;
      dct_coeffs[19][29] = 32'h00C8FB2F;
      dct_coeffs[19][30] = 32'h0F109082;
      dct_coeffs[19][31] = 32'hF6780402;
      dct_coeffs[20][0] = 32'h08E39D9C;
      dct_coeffs[20][1] = 32'hF04EB419;
      dct_coeffs[20][2] = 32'h031F1707;
      dct_coeffs[20][3] = 32'h0D4DB314;
      dct_coeffs[20][4] = 32'hF2B24CEC;
      dct_coeffs[20][5] = 32'hFCE0E8F9;
      dct_coeffs[20][6] = 32'h0FB14BE7;
      dct_coeffs[20][7] = 32'hF71C6264;
      dct_coeffs[20][8] = 32'hF71C6264;
      dct_coeffs[20][9] = 32'h0FB14BE7;
      dct_coeffs[20][10] = 32'hFCE0E8F9;
      dct_coeffs[20][11] = 32'hF2B24CEC;
      dct_coeffs[20][12] = 32'h0D4DB314;
      dct_coeffs[20][13] = 32'h031F1707;
      dct_coeffs[20][14] = 32'hF04EB419;
      dct_coeffs[20][15] = 32'h08E39D9C;
      dct_coeffs[20][16] = 32'h08E39D9C;
      dct_coeffs[20][17] = 32'hF04EB419;
      dct_coeffs[20][18] = 32'h031F1707;
      dct_coeffs[20][19] = 32'h0D4DB314;
      dct_coeffs[20][20] = 32'hF2B24CEC;
      dct_coeffs[20][21] = 32'hFCE0E8F9;
      dct_coeffs[20][22] = 32'h0FB14BE7;
      dct_coeffs[20][23] = 32'hF71C6264;
      dct_coeffs[20][24] = 32'hF71C6264;
      dct_coeffs[20][25] = 32'h0FB14BE7;
      dct_coeffs[20][26] = 32'hFCE0E8F9;
      dct_coeffs[20][27] = 32'hF2B24CEC;
      dct_coeffs[20][28] = 32'h0D4DB314;
      dct_coeffs[20][29] = 32'h031F1707;
      dct_coeffs[20][30] = 32'hF04EB419;
      dct_coeffs[20][31] = 32'h08E39D9C;
      dct_coeffs[21][0] = 32'h0839C3CC;
      dct_coeffs[21][1] = 32'hF004EF0F;
      dct_coeffs[21][2] = 32'h06D74402;
      dct_coeffs[21][3] = 32'h0987FBFE;
      dct_coeffs[21][4] = 32'hF02C5541;
      dct_coeffs[21][5] = 32'h0563E69D;
      dct_coeffs[21][6] = 32'h0ABEB49A;
      dct_coeffs[21][7] = 32'hF07AC083;
      dct_coeffs[21][8] = 32'h03E33F2F;
      dct_coeffs[21][9] = 32'h0BDAEF91;
      dct_coeffs[21][10] = 32'hF0EF6F7E;
      dct_coeffs[21][11] = 32'h0259020D;
      dct_coeffs[21][12] = 32'h0CD9F023;
      dct_coeffs[21][13] = 32'hF1894286;
      dct_coeffs[21][14] = 32'h00C8FB2F;
      dct_coeffs[21][15] = 32'h0DB941A2;
      dct_coeffs[21][16] = 32'hF246BE5E;
      dct_coeffs[21][17] = 32'hFF3704D1;
      dct_coeffs[21][18] = 32'h0E76BD7A;
      dct_coeffs[21][19] = 32'hF3260FDD;
      dct_coeffs[21][20] = 32'hFDA6FDF3;
      dct_coeffs[21][21] = 32'h0F109082;
      dct_coeffs[21][22] = 32'hF425106F;
      dct_coeffs[21][23] = 32'hFC1CC0D1;
      dct_coeffs[21][24] = 32'h0F853F7D;
      dct_coeffs[21][25] = 32'hF5414B66;
      dct_coeffs[21][26] = 32'hFA9C1963;
      dct_coeffs[21][27] = 32'h0FD3AABF;
      dct_coeffs[21][28] = 32'hF6780402;
      dct_coeffs[21][29] = 32'hF928BBFE;
      dct_coeffs[21][30] = 32'h0FFB10F1;
      dct_coeffs[21][31] = 32'hF7C63C34;
      dct_coeffs[22][0] = 32'h078AD74E;
      dct_coeffs[22][1] = 32'hF013B92F;
      dct_coeffs[22][2] = 32'h0A267992;
      dct_coeffs[22][3] = 32'h04A5018B;
      dct_coeffs[22][4] = 32'hF0B05F55;
      dct_coeffs[22][5] = 32'h0C5E4035;
      dct_coeffs[22][6] = 32'h01917A6B;
      dct_coeffs[22][7] = 32'hF1E3A688;
      dct_coeffs[22][8] = 32'h0E1C5978;
      dct_coeffs[22][9] = 32'hFE6E8595;
      dct_coeffs[22][10] = 32'hF3A1BFCB;
      dct_coeffs[22][11] = 32'h0F4FA0AB;
      dct_coeffs[22][12] = 32'hFB5AFE75;
      dct_coeffs[22][13] = 32'hF5D9866E;
      dct_coeffs[22][14] = 32'h0FEC46D1;
      dct_coeffs[22][15] = 32'hF87528B2;
      dct_coeffs[22][16] = 32'hF87528B2;
      dct_coeffs[22][17] = 32'h0FEC46D1;
      dct_coeffs[22][18] = 32'hF5D9866E;
      dct_coeffs[22][19] = 32'hFB5AFE75;
      dct_coeffs[22][20] = 32'h0F4FA0AB;
      dct_coeffs[22][21] = 32'hF3A1BFCB;
      dct_coeffs[22][22] = 32'hFE6E8595;
      dct_coeffs[22][23] = 32'h0E1C5978;
      dct_coeffs[22][24] = 32'hF1E3A688;
      dct_coeffs[22][25] = 32'h01917A6B;
      dct_coeffs[22][26] = 32'h0C5E4035;
      dct_coeffs[22][27] = 32'hF0B05F55;
      dct_coeffs[22][28] = 32'h04A5018B;
      dct_coeffs[22][29] = 32'h0A267992;
      dct_coeffs[22][30] = 32'hF013B92F;
      dct_coeffs[22][31] = 32'h078AD74E;
      dct_coeffs[23][0] = 32'h06D74402;
      dct_coeffs[23][1] = 32'hF07AC083;
      dct_coeffs[23][2] = 32'h0CD9F023;
      dct_coeffs[23][3] = 32'hFF3704D1;
      dct_coeffs[23][4] = 32'hF425106F;
      dct_coeffs[23][5] = 32'h0FD3AABF;
      dct_coeffs[23][6] = 32'hF7C63C34;
      dct_coeffs[23][7] = 32'hFA9C1963;
      dct_coeffs[23][8] = 32'h0F109082;
      dct_coeffs[23][9] = 32'hF246BE5E;
      dct_coeffs[23][10] = 32'h0259020D;
      dct_coeffs[23][11] = 32'h0ABEB49A;
      dct_coeffs[23][12] = 32'hF004EF0F;
      dct_coeffs[23][13] = 32'h0987FBFE;
      dct_coeffs[23][14] = 32'h03E33F2F;
      dct_coeffs[23][15] = 32'hF1894286;
      dct_coeffs[23][16] = 32'h0E76BD7A;
      dct_coeffs[23][17] = 32'hFC1CC0D1;
      dct_coeffs[23][18] = 32'hF6780402;
      dct_coeffs[23][19] = 32'h0FFB10F1;
      dct_coeffs[23][20] = 32'hF5414B66;
      dct_coeffs[23][21] = 32'hFDA6FDF3;
      dct_coeffs[23][22] = 32'h0DB941A2;
      dct_coeffs[23][23] = 32'hF0EF6F7E;
      dct_coeffs[23][24] = 32'h0563E69D;
      dct_coeffs[23][25] = 32'h0839C3CC;
      dct_coeffs[23][26] = 32'hF02C5541;
      dct_coeffs[23][27] = 32'h0BDAEF91;
      dct_coeffs[23][28] = 32'h00C8FB2F;
      dct_coeffs[23][29] = 32'hF3260FDD;
      dct_coeffs[23][30] = 32'h0F853F7D;
      dct_coeffs[23][31] = 32'hF928BBFE;
      dct_coeffs[24][0] = 32'h061F78A9;
      dct_coeffs[24][1] = 32'hF137CA19;
      dct_coeffs[24][2] = 32'h0EC835E7;
      dct_coeffs[24][3] = 32'hF9E08757;
      dct_coeffs[24][4] = 32'hF9E08757;
      dct_coeffs[24][5] = 32'h0EC835E7;
      dct_coeffs[24][6] = 32'hF137CA19;
      dct_coeffs[24][7] = 32'h061F78A9;
      dct_coeffs[24][8] = 32'h061F78A9;
      dct_coeffs[24][9] = 32'hF137CA19;
      dct_coeffs[24][10] = 32'h0EC835E7;
      dct_coeffs[24][11] = 32'hF9E08757;
      dct_coeffs[24][12] = 32'hF9E08757;
      dct_coeffs[24][13] = 32'h0EC835E7;
      dct_coeffs[24][14] = 32'hF137CA19;
      dct_coeffs[24][15] = 32'h061F78A9;
      dct_coeffs[24][16] = 32'h061F78A9;
      dct_coeffs[24][17] = 32'hF137CA19;
      dct_coeffs[24][18] = 32'h0EC835E7;
      dct_coeffs[24][19] = 32'hF9E08757;
      dct_coeffs[24][20] = 32'hF9E08757;
      dct_coeffs[24][21] = 32'h0EC835E7;
      dct_coeffs[24][22] = 32'hF137CA19;
      dct_coeffs[24][23] = 32'h061F78A9;
      dct_coeffs[24][24] = 32'h061F78A9;
      dct_coeffs[24][25] = 32'hF137CA19;
      dct_coeffs[24][26] = 32'h0EC835E7;
      dct_coeffs[24][27] = 32'hF9E08757;
      dct_coeffs[24][28] = 32'hF9E08757;
      dct_coeffs[24][29] = 32'h0EC835E7;
      dct_coeffs[24][30] = 32'hF137CA19;
      dct_coeffs[24][31] = 32'h061F78A9;
      dct_coeffs[25][0] = 32'h0563E69D;
      dct_coeffs[25][1] = 32'hF246BE5E;
      dct_coeffs[25][2] = 32'h0FD3AABF;
      dct_coeffs[25][3] = 32'hF5414B66;
      dct_coeffs[25][4] = 32'h00C8FB2F;
      dct_coeffs[25][5] = 32'h0987FBFE;
      dct_coeffs[25][6] = 32'hF07AC083;
      dct_coeffs[25][7] = 32'h0E76BD7A;
      dct_coeffs[25][8] = 32'hF928BBFE;
      dct_coeffs[25][9] = 32'hFC1CC0D1;
      dct_coeffs[25][10] = 32'h0CD9F023;
      dct_coeffs[25][11] = 32'hF004EF0F;
      dct_coeffs[25][12] = 32'h0BDAEF91;
      dct_coeffs[25][13] = 32'hFDA6FDF3;
      dct_coeffs[25][14] = 32'hF7C63C34;
      dct_coeffs[25][15] = 32'h0F109082;
      dct_coeffs[25][16] = 32'hF0EF6F7E;
      dct_coeffs[25][17] = 32'h0839C3CC;
      dct_coeffs[25][18] = 32'h0259020D;
      dct_coeffs[25][19] = 32'hF425106F;
      dct_coeffs[25][20] = 32'h0FFB10F1;
      dct_coeffs[25][21] = 32'hF3260FDD;
      dct_coeffs[25][22] = 32'h03E33F2F;
      dct_coeffs[25][23] = 32'h06D74402;
      dct_coeffs[25][24] = 32'hF1894286;
      dct_coeffs[25][25] = 32'h0F853F7D;
      dct_coeffs[25][26] = 32'hF6780402;
      dct_coeffs[25][27] = 32'hFF3704D1;
      dct_coeffs[25][28] = 32'h0ABEB49A;
      dct_coeffs[25][29] = 32'hF02C5541;
      dct_coeffs[25][30] = 32'h0DB941A2;
      dct_coeffs[25][31] = 32'hFA9C1963;
      dct_coeffs[26][0] = 32'h04A5018B;
      dct_coeffs[26][1] = 32'hF3A1BFCB;
      dct_coeffs[26][2] = 32'h0FEC46D1;
      dct_coeffs[26][3] = 32'hF1E3A688;
      dct_coeffs[26][4] = 32'h078AD74E;
      dct_coeffs[26][5] = 32'h01917A6B;
      dct_coeffs[26][6] = 32'hF5D9866E;
      dct_coeffs[26][7] = 32'h0F4FA0AB;
      dct_coeffs[26][8] = 32'hF0B05F55;
      dct_coeffs[26][9] = 32'h0A267992;
      dct_coeffs[26][10] = 32'hFE6E8595;
      dct_coeffs[26][11] = 32'hF87528B2;
      dct_coeffs[26][12] = 32'h0E1C5978;
      dct_coeffs[26][13] = 32'hF013B92F;
      dct_coeffs[26][14] = 32'h0C5E4035;
      dct_coeffs[26][15] = 32'hFB5AFE75;
      dct_coeffs[26][16] = 32'hFB5AFE75;
      dct_coeffs[26][17] = 32'h0C5E4035;
      dct_coeffs[26][18] = 32'hF013B92F;
      dct_coeffs[26][19] = 32'h0E1C5978;
      dct_coeffs[26][20] = 32'hF87528B2;
      dct_coeffs[26][21] = 32'hFE6E8595;
      dct_coeffs[26][22] = 32'h0A267992;
      dct_coeffs[26][23] = 32'hF0B05F55;
      dct_coeffs[26][24] = 32'h0F4FA0AB;
      dct_coeffs[26][25] = 32'hF5D9866E;
      dct_coeffs[26][26] = 32'h01917A6B;
      dct_coeffs[26][27] = 32'h078AD74E;
      dct_coeffs[26][28] = 32'hF1E3A688;
      dct_coeffs[26][29] = 32'h0FEC46D1;
      dct_coeffs[26][30] = 32'hF3A1BFCB;
      dct_coeffs[26][31] = 32'h04A5018B;
      dct_coeffs[27][0] = 32'h03E33F2F;
      dct_coeffs[27][1] = 32'hF5414B66;
      dct_coeffs[27][2] = 32'h0F109082;
      dct_coeffs[27][3] = 32'hF02C5541;
      dct_coeffs[27][4] = 32'h0CD9F023;
      dct_coeffs[27][5] = 32'hF928BBFE;
      dct_coeffs[27][6] = 32'hFF3704D1;
      dct_coeffs[27][7] = 32'h0839C3CC;
      dct_coeffs[27][8] = 32'hF246BE5E;
      dct_coeffs[27][9] = 32'h0FFB10F1;
      dct_coeffs[27][10] = 32'hF1894286;
      dct_coeffs[27][11] = 32'h0987FBFE;
      dct_coeffs[27][12] = 32'hFDA6FDF3;
      dct_coeffs[27][13] = 32'hFA9C1963;
      dct_coeffs[27][14] = 32'h0BDAEF91;
      dct_coeffs[27][15] = 32'hF07AC083;
      dct_coeffs[27][16] = 32'h0F853F7D;
      dct_coeffs[27][17] = 32'hF425106F;
      dct_coeffs[27][18] = 32'h0563E69D;
      dct_coeffs[27][19] = 32'h0259020D;
      dct_coeffs[27][20] = 32'hF6780402;
      dct_coeffs[27][21] = 32'h0E76BD7A;
      dct_coeffs[27][22] = 32'hF004EF0F;
      dct_coeffs[27][23] = 32'h0DB941A2;
      dct_coeffs[27][24] = 32'hF7C63C34;
      dct_coeffs[27][25] = 32'h00C8FB2F;
      dct_coeffs[27][26] = 32'h06D74402;
      dct_coeffs[27][27] = 32'hF3260FDD;
      dct_coeffs[27][28] = 32'h0FD3AABF;
      dct_coeffs[27][29] = 32'hF0EF6F7E;
      dct_coeffs[27][30] = 32'h0ABEB49A;
      dct_coeffs[27][31] = 32'hFC1CC0D1;
      dct_coeffs[28][0] = 32'h031F1707;
      dct_coeffs[28][1] = 32'hF71C6264;
      dct_coeffs[28][2] = 32'h0D4DB314;
      dct_coeffs[28][3] = 32'hF04EB419;
      dct_coeffs[28][4] = 32'h0FB14BE7;
      dct_coeffs[28][5] = 32'hF2B24CEC;
      dct_coeffs[28][6] = 32'h08E39D9C;
      dct_coeffs[28][7] = 32'hFCE0E8F9;
      dct_coeffs[28][8] = 32'hFCE0E8F9;
      dct_coeffs[28][9] = 32'h08E39D9C;
      dct_coeffs[28][10] = 32'hF2B24CEC;
      dct_coeffs[28][11] = 32'h0FB14BE7;
      dct_coeffs[28][12] = 32'hF04EB419;
      dct_coeffs[28][13] = 32'h0D4DB314;
      dct_coeffs[28][14] = 32'hF71C6264;
      dct_coeffs[28][15] = 32'h031F1707;
      dct_coeffs[28][16] = 32'h031F1707;
      dct_coeffs[28][17] = 32'hF71C6264;
      dct_coeffs[28][18] = 32'h0D4DB314;
      dct_coeffs[28][19] = 32'hF04EB419;
      dct_coeffs[28][20] = 32'h0FB14BE7;
      dct_coeffs[28][21] = 32'hF2B24CEC;
      dct_coeffs[28][22] = 32'h08E39D9C;
      dct_coeffs[28][23] = 32'hFCE0E8F9;
      dct_coeffs[28][24] = 32'hFCE0E8F9;
      dct_coeffs[28][25] = 32'h08E39D9C;
      dct_coeffs[28][26] = 32'hF2B24CEC;
      dct_coeffs[28][27] = 32'h0FB14BE7;
      dct_coeffs[28][28] = 32'hF04EB419;
      dct_coeffs[28][29] = 32'h0D4DB314;
      dct_coeffs[28][30] = 32'hF71C6264;
      dct_coeffs[28][31] = 32'h031F1707;
      dct_coeffs[29][0] = 32'h0259020D;
      dct_coeffs[29][1] = 32'hF928BBFE;
      dct_coeffs[29][2] = 32'h0ABEB49A;
      dct_coeffs[29][3] = 32'hF246BE5E;
      dct_coeffs[29][4] = 32'h0F853F7D;
      dct_coeffs[29][5] = 32'hF004EF0F;
      dct_coeffs[29][6] = 32'h0F109082;
      dct_coeffs[29][7] = 32'hF3260FDD;
      dct_coeffs[29][8] = 32'h0987FBFE;
      dct_coeffs[29][9] = 32'hFA9C1963;
      dct_coeffs[29][10] = 32'h00C8FB2F;
      dct_coeffs[29][11] = 32'h03E33F2F;
      dct_coeffs[29][12] = 32'hF7C63C34;
      dct_coeffs[29][13] = 32'h0BDAEF91;
      dct_coeffs[29][14] = 32'hF1894286;
      dct_coeffs[29][15] = 32'h0FD3AABF;
      dct_coeffs[29][16] = 32'hF02C5541;
      dct_coeffs[29][17] = 32'h0E76BD7A;
      dct_coeffs[29][18] = 32'hF425106F;
      dct_coeffs[29][19] = 32'h0839C3CC;
      dct_coeffs[29][20] = 32'hFC1CC0D1;
      dct_coeffs[29][21] = 32'hFF3704D1;
      dct_coeffs[29][22] = 32'h0563E69D;
      dct_coeffs[29][23] = 32'hF6780402;
      dct_coeffs[29][24] = 32'h0CD9F023;
      dct_coeffs[29][25] = 32'hF0EF6F7E;
      dct_coeffs[29][26] = 32'h0FFB10F1;
      dct_coeffs[29][27] = 32'hF07AC083;
      dct_coeffs[29][28] = 32'h0DB941A2;
      dct_coeffs[29][29] = 32'hF5414B66;
      dct_coeffs[29][30] = 32'h06D74402;
      dct_coeffs[29][31] = 32'hFDA6FDF3;
      dct_coeffs[30][0] = 32'h01917A6B;
      dct_coeffs[30][1] = 32'hFB5AFE75;
      dct_coeffs[30][2] = 32'h078AD74E;
      dct_coeffs[30][3] = 32'hF5D9866E;
      dct_coeffs[30][4] = 32'h0C5E4035;
      dct_coeffs[30][5] = 32'hF1E3A688;
      dct_coeffs[30][6] = 32'h0F4FA0AB;
      dct_coeffs[30][7] = 32'hF013B92F;
      dct_coeffs[30][8] = 32'h0FEC46D1;
      dct_coeffs[30][9] = 32'hF0B05F55;
      dct_coeffs[30][10] = 32'h0E1C5978;
      dct_coeffs[30][11] = 32'hF3A1BFCB;
      dct_coeffs[30][12] = 32'h0A267992;
      dct_coeffs[30][13] = 32'hF87528B2;
      dct_coeffs[30][14] = 32'h04A5018B;
      dct_coeffs[30][15] = 32'hFE6E8595;
      dct_coeffs[30][16] = 32'hFE6E8595;
      dct_coeffs[30][17] = 32'h04A5018B;
      dct_coeffs[30][18] = 32'hF87528B2;
      dct_coeffs[30][19] = 32'h0A267992;
      dct_coeffs[30][20] = 32'hF3A1BFCB;
      dct_coeffs[30][21] = 32'h0E1C5978;
      dct_coeffs[30][22] = 32'hF0B05F55;
      dct_coeffs[30][23] = 32'h0FEC46D1;
      dct_coeffs[30][24] = 32'hF013B92F;
      dct_coeffs[30][25] = 32'h0F4FA0AB;
      dct_coeffs[30][26] = 32'hF1E3A688;
      dct_coeffs[30][27] = 32'h0C5E4035;
      dct_coeffs[30][28] = 32'hF5D9866E;
      dct_coeffs[30][29] = 32'h078AD74E;
      dct_coeffs[30][30] = 32'hFB5AFE75;
      dct_coeffs[30][31] = 32'h01917A6B;
      dct_coeffs[31][0] = 32'h00C8FB2F;
      dct_coeffs[31][1] = 32'hFDA6FDF3;
      dct_coeffs[31][2] = 32'h03E33F2F;
      dct_coeffs[31][3] = 32'hFA9C1963;
      dct_coeffs[31][4] = 32'h06D74402;
      dct_coeffs[31][5] = 32'hF7C63C34;
      dct_coeffs[31][6] = 32'h0987FBFE;
      dct_coeffs[31][7] = 32'hF5414B66;
      dct_coeffs[31][8] = 32'h0BDAEF91;
      dct_coeffs[31][9] = 32'hF3260FDD;
      dct_coeffs[31][10] = 32'h0DB941A2;
      dct_coeffs[31][11] = 32'hF1894286;
      dct_coeffs[31][12] = 32'h0F109082;
      dct_coeffs[31][13] = 32'hF07AC083;
      dct_coeffs[31][14] = 32'h0FD3AABF;
      dct_coeffs[31][15] = 32'hF004EF0F;
      dct_coeffs[31][16] = 32'h0FFB10F1;
      dct_coeffs[31][17] = 32'hF02C5541;
      dct_coeffs[31][18] = 32'h0F853F7D;
      dct_coeffs[31][19] = 32'hF0EF6F7E;
      dct_coeffs[31][20] = 32'h0E76BD7A;
      dct_coeffs[31][21] = 32'hF246BE5E;
      dct_coeffs[31][22] = 32'h0CD9F023;
      dct_coeffs[31][23] = 32'hF425106F;
      dct_coeffs[31][24] = 32'h0ABEB49A;
      dct_coeffs[31][25] = 32'hF6780402;
      dct_coeffs[31][26] = 32'h0839C3CC;
      dct_coeffs[31][27] = 32'hF928BBFE;
      dct_coeffs[31][28] = 32'h0563E69D;
      dct_coeffs[31][29] = 32'hFC1CC0D1;
      dct_coeffs[31][30] = 32'h0259020D;
      dct_coeffs[31][31] = 32'hFF3704D1;

end

endmodule
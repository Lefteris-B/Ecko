module dct_module #(
  parameter Q_L = 11,  // Number of fractional bits for logarithm output
  parameter Q_D = 4,   // Number of fractional bits for DCT output
  parameter N = 32     // Size of the DCT input vector
) (
  input wire clk,
  input wire rst,
  input wire signed [Q_L-1:0] data_in,
  input wire data_valid,
  output reg signed [Q_D-1:0] dct_out,
  output reg dct_valid
);

  localparam COEFF_WIDTH = 16;

  reg signed [Q_L-1:0] input_buffer [0:N-1];
  reg [$clog2(N)-1:0] input_counter;
  reg [$clog2(N)-1:0] output_counter;
  reg signed [COEFF_WIDTH-1:0] coeff;
  reg signed [Q_L+COEFF_WIDTH-1:0] mult;
  reg signed [Q_L+COEFF_WIDTH-1:0] accumulator;
  reg [1:0] state;

  // Precomputed fixed-point DCT coefficients (Chen's algorithm for N=32)
  always @(*) begin
    case (output_counter)
     0: coeff = (input_counter == 0) ? 0x16a1 : (input_counter == 1) ? 0x16a1 : (input_counter == 2) ? 0x16a1 : (input_counter == 3) ? 0x16a1 : (input_counter == 4) ? 0x16a1 : (input_counter == 5) ? 0x16a1 : (input_counter == 6) ? 0x16a1 : (input_counter == 7) ? 0x16a1 : (input_counter == 8) ? 0x16a1 : (input_counter == 9) ? 0x16a1 : (input_counter == 10) ? 0x16a1 : (input_counter == 11) ? 0x16a1 : (input_counter == 12) ? 0x16a1 : (input_counter == 13) ? 0x16a1 : (input_counter == 14) ? 0x16a1 : (input_counter == 15) ? 0x16a1 : (input_counter == 16) ? 0x16a1 : (input_counter == 17) ? 0x16a1 : (input_counter == 18) ? 0x16a1 : (input_counter == 19) ? 0x16a1 : (input_counter == 20) ? 0x16a1 : (input_counter == 21) ? 0x16a1 : (input_counter == 22) ? 0x16a1 : (input_counter == 23) ? 0x16a1 : (input_counter == 24) ? 0x16a1 : (input_counter == 25) ? 0x16a1 : (input_counter == 26) ? 0x16a1 : (input_counter == 27) ? 0x16a1 : (input_counter == 28) ? 0x16a1 : (input_counter == 29) ? 0x16a1 : (input_counter == 30) ? 0x16a1 : 0x16a1;
1: coeff = (input_counter == 0) ? 0x1ff6 : (input_counter == 1) ? 0x1fa7 : (input_counter == 2) ? 0x1f0a : (input_counter == 3) ? 0x1e21 : (input_counter == 4) ? 0x1ced : (input_counter == 5) ? 0x1b73 : (input_counter == 6) ? 0x19b4 : (input_counter == 7) ? 0x17b6 : (input_counter == 8) ? 0x157d : (input_counter == 9) ? 0x1310 : (input_counter == 10) ? 0x1074 : (input_counter == 11) ? 0x0daf : (input_counter == 12) ? 0x0ac8 : (input_counter == 13) ? 0x07c6 : (input_counter == 14) ? 0x04b2 : (input_counter == 15) ? 0x0192 : (input_counter == 16) ? -0x192 : (input_counter == 17) ? -0x4b2 : (input_counter == 18) ? -0x7c6 : (input_counter == 19) ? -0xac8 : (input_counter == 20) ? -0xdaf : (input_counter == 21) ? -0x1074 : (input_counter == 22) ? -0x1310 : (input_counter == 23) ? -0x157d : (input_counter == 24) ? -0x17b6 : (input_counter == 25) ? -0x19b4 : (input_counter == 26) ? -0x1b73 : (input_counter == 27) ? -0x1ced : (input_counter == 28) ? -0x1e21 : (input_counter == 29) ? -0x1f0a : (input_counter == 30) ? -0x1fa7 : -0x1ff6;
2: coeff = (input_counter == 0) ? 0x1fd9 : (input_counter == 1) ? 0x1e9f : (input_counter == 2) ? 0x1c39 : (input_counter == 3) ? 0x18bd : (input_counter == 4) ? 0x144d : (input_counter == 5) ? 0x0f16 : (input_counter == 6) ? 0x094a : (input_counter == 7) ? 0x0323 : (input_counter == 8) ? -0x323 : (input_counter == 9) ? -0x94a : (input_counter == 10) ? -0xf16 : (input_counter == 11) ? -0x144d : (input_counter == 12) ? -0x18bd : (input_counter == 13) ? -0x1c39 : (input_counter == 14) ? -0x1e9f : (input_counter == 15) ? -0x1fd9 : (input_counter == 16) ? -0x1fd9 : (input_counter == 17) ? -0x1e9f : (input_counter == 18) ? -0x1c39 : (input_counter == 19) ? -0x18bd : (input_counter == 20) ? -0x144d : (input_counter == 21) ? -0xf16 : (input_counter == 22) ? -0x94a : (input_counter == 23) ? -0x323 : (input_counter == 24) ? 0x0323 : (input_counter == 25) ? 0x094a : (input_counter == 26) ? 0x0f16 : (input_counter == 27) ? 0x144d : (input_counter == 28) ? 0x18bd : (input_counter == 29) ? 0x1c39 : (input_counter == 30) ? 0x1e9f : 0x1fd9;
3: coeff = (input_counter == 0) ? 0x1fa7 : (input_counter == 1) ? 0x1ced : (input_counter == 2) ? 0x17b6 : (input_counter == 3) ? 0x1074 : (input_counter == 4) ? 0x07c6 : (input_counter == 5) ? -0x192 : (input_counter == 6) ? -0xac8 : (input_counter == 7) ? -0x1310 : (input_counter == 8) ? -0x19b4 : (input_counter == 9) ? -0x1e21 : (input_counter == 10) ? -0x1ff6 : (input_counter == 11) ? -0x1f0a : (input_counter == 12) ? -0x1b73 : (input_counter == 13) ? -0x157d : (input_counter == 14) ? -0xdaf : (input_counter == 15) ? -0x4b2 : (input_counter == 16) ? 0x04b2 : (input_counter == 17) ? 0x0daf : (input_counter == 18) ? 0x157d : (input_counter == 19) ? 0x1b73 : (input_counter == 20) ? 0x1f0a : (input_counter == 21) ? 0x1ff6 : (input_counter == 22) ? 0x1e21 : (input_counter == 23) ? 0x19b4 : (input_counter == 24) ? 0x1310 : (input_counter == 25) ? 0x0ac8 : (input_counter == 26) ? 0x0192 : (input_counter == 27) ? -0x7c6 : (input_counter == 28) ? -0x1074 : (input_counter == 29) ? -0x17b6 : (input_counter == 30) ? -0x1ced : -0x1fa7;
4: coeff = (input_counter == 0) ? 0x1f63 : (input_counter == 1) ? 0x1a9b : (input_counter == 2) ? 0x11c7 : (input_counter == 3) ? 0x063e : (input_counter == 4) ? -0x63e : (input_counter == 5) ? -0x11c7 : (input_counter == 6) ? -0x1a9b : (input_counter == 7) ? -0x1f63 : (input_counter == 8) ? -0x1f63 : (input_counter == 9) ? -0x1a9b : (input_counter == 10) ? -0x11c7 : (input_counter == 11) ? -0x63e : (input_counter == 12) ? 0x063e : (input_counter == 13) ? 0x11c7 : (input_counter == 14) ? 0x1a9b : (input_counter == 15) ? 0x1f63 : (input_counter == 16) ? 0x1f63 : (input_counter == 17) ? 0x1a9b : (input_counter == 18) ? 0x11c7 : (input_counter == 19) ? 0x063e : (input_counter == 20) ? -0x63e : (input_counter == 21) ? -0x11c7 : (input_counter == 22) ? -0x1a9b : (input_counter == 23) ? -0x1f63 : (input_counter == 24) ? -0x1f63 : (input_counter == 25) ? -0x1a9b : (input_counter == 26) ? -0x11c7 : (input_counter == 27) ? -0x63e : (input_counter == 28) ? 0x063e : (input_counter == 29) ? 0x11c7 : (input_counter == 30) ? 0x1a9b : 0x1f63;
5: coeff = (input_counter == 0) ? 0x1f0a : (input_counter == 1) ? 0x17b6 : (input_counter == 2) ? 0x0ac8 : (input_counter == 3) ? -0x4b2 : (input_counter == 4) ? -0x1310 : (input_counter == 5) ? -0x1ced : (input_counter == 6) ? -0x1ff6 : (input_counter == 7) ? -0x1b73 : (input_counter == 8) ? -0x1074 : (input_counter == 9) ? -0x192 : (input_counter == 10) ? 0x0daf : (input_counter == 11) ? 0x19b4 : (input_counter == 12) ? 0x1fa7 : (input_counter == 13) ? 0x1e21 : (input_counter == 14) ? 0x157d : (input_counter == 15) ? 0x07c6 : (input_counter == 16) ? -0x7c6 : (input_counter == 17) ? -0x157d : (input_counter == 18) ? -0x1e21 : (input_counter == 19) ? -0x1fa7 : (input_counter == 20) ? -0x19b4 : (input_counter == 21) ? -0xdaf : (input_counter == 22) ? 0x0192 : (input_counter == 23) ? 0x1074 : (input_counter == 24) ? 0x1b73 : (input_counter == 25) ? 0x1ff6 : (input_counter == 26) ? 0x1ced : (input_counter == 27) ? 0x1310 : (input_counter == 28) ? 0x04b2 : (input_counter == 29) ? -0xac8 : (input_counter == 30) ? -0x17b6 : -0x1f0a;
6: coeff = (input_counter == 0) ? 0x1e9f : (input_counter == 1) ? 0x144d : (input_counter == 2) ? 0x0323 : (input_counter == 3) ? -0xf16 : (input_counter == 4) ? -0x1c39 : (input_counter == 5) ? -0x1fd9 : (input_counter == 6) ? -0x18bd : (input_counter == 7) ? -0x94a : (input_counter == 8) ? 0x094a : (input_counter == 9) ? 0x18bd : (input_counter == 10) ? 0x1fd9 : (input_counter == 11) ? 0x1c39 : (input_counter == 12) ? 0x0f16 : (input_counter == 13) ? -0x323 : (input_counter == 14) ? -0x144d : (input_counter == 15) ? -0x1e9f : (input_counter == 16) ? -0x1e9f : (input_counter == 17) ? -0x144d : (input_counter == 18) ? -0x323 : (input_counter == 19) ? 0x0f16 : (input_counter == 20) ? 0x1c39 : (input_counter == 21) ? 0x1fd9 : (input_counter == 22) ? 0x18bd : (input_counter == 23) ? 0x094a : (input_counter == 24) ? -0x94a : (input_counter == 25) ? -0x18bd : (input_counter == 26) ? -0x1fd9 : (input_counter == 27) ? -0x1c39 : (input_counter == 28) ? -0xf16 : (input_counter == 29) ? 0x0323 : (input_counter == 30) ? 0x144d : 0x1e9f;
7: coeff = (input_counter == 0) ? 0x1e21 : (input_counter == 1) ? 0x1074 : (input_counter == 2) ? -0x4b2 : (input_counter == 3) ? -0x17b6 : (input_counter == 4) ? -0x1ff6 : (input_counter == 5) ? -0x19b4 : (input_counter == 6) ? -0x7c6 : (input_counter == 7) ? 0x0daf : (input_counter == 8) ? 0x1ced : (input_counter == 9) ? 0x1f0a : (input_counter == 10) ? 0x1310 : (input_counter == 11) ? -0x192 : (input_counter == 12) ? -0x157d : (input_counter == 13) ? -0x1fa7 : (input_counter == 14) ? -0x1b73 : (input_counter == 15) ? -0xac8 : (input_counter == 16) ? 0x0ac8 : (input_counter == 17) ? 0x1b73 : (input_counter == 18) ? 0x1fa7 : (input_counter == 19) ? 0x157d : (input_counter == 20) ? 0x0192 : (input_counter == 21) ? -0x1310 : (input_counter == 22) ? -0x1f0a : (input_counter == 23) ? -0x1ced : (input_counter == 24) ? -0xdaf : (input_counter == 25) ? 0x07c6 : (input_counter == 26) ? 0x19b4 : (input_counter == 27) ? 0x1ff6 : (input_counter == 28) ? 0x17b6 : (input_counter == 29) ? 0x04b2 : (input_counter == 30) ? -0x1074 : -0x1e21;
8: coeff = (input_counter == 0) ? 0x1d90 : (input_counter == 1) ? 0x0c3f : (input_counter == 2) ? -0xc3f : (input_counter == 3) ? -0x1d90 : (input_counter == 4) ? -0x1d90 : (input_counter == 5) ? -0xc3f : (input_counter == 6) ? 0x0c3f : (input_counter == 7) ? 0x1d90 : (input_counter == 8) ? 0x1d90 : (input_counter == 9) ? 0x0c3f : (input_counter == 10) ? -0xc3f : (input_counter == 11) ? -0x1d90 : (input_counter == 12) ? -0x1d90 : (input_counter == 13) ? -0xc3f : (input_counter == 14) ? 0x0c3f : (input_counter == 15) ? 0x1d90 : (input_counter == 16) ? 0x1d90 : (input_counter == 17) ? 0x0c3f : (input_counter == 18) ? -0xc3f : (input_counter == 19) ? -0x1d90 : (input_counter == 20) ? -0x1d90 : (input_counter == 21) ? -0xc3f : (input_counter == 22) ? 0x0c3f : (input_counter == 23) ? 0x1d90 : (input_counter == 24) ? 0x1d90 : (input_counter == 25) ? 0x0c3f : (input_counter == 26) ? -0xc3f : (input_counter == 27) ? -0x1d90 : (input_counter == 28) ? -0x1d90 : (input_counter == 29) ? -0xc3f : (input_counter == 30) ? 0x0c3f : 0x1d90;
9: coeff = (input_counter == 0) ? 0x1ced : (input_counter == 1) ? 0x07c6 : (input_counter == 2) ? -0x1310 : (input_counter == 3) ? -0x1ff6 : (input_counter == 4) ? -0x157d : (input_counter == 5) ? 0x04b2 : (input_counter == 6) ? 0x1b73 : (input_counter == 7) ? 0x1e21 : (input_counter == 8) ? 0x0ac8 : (input_counter == 9) ? -0x1074 : (input_counter == 10) ? -0x1fa7 : (input_counter == 11) ? -0x17b6 : (input_counter == 12) ? 0x0192 : (input_counter == 13) ? 0x19b4 : (input_counter == 14) ? 0x1f0a : (input_counter == 15) ? 0x0daf : (input_counter == 16) ? -0xdaf : (input_counter == 17) ? -0x1f0a : (input_counter == 18) ? -0x19b4 : (input_counter == 19) ? -0x192 : (input_counter == 20) ? 0x17b6 : (input_counter == 21) ? 0x1fa7 : (input_counter == 22) ? 0x1074 : (input_counter == 23) ? -0xac8 : (input_counter == 24) ? -0x1e21 : (input_counter == 25) ? -0x1b73 : (input_counter == 26) ? -0x4b2 : (input_counter == 27) ? 0x157d : (input_counter == 28) ? 0x1ff6 : (input_counter == 29) ? 0x1310 : (input_counter == 30) ? -0x7c6 : -0x1ced;
10: coeff = (input_counter == 0) ? 0x1c39 : (input_counter == 1) ? 0x0323 : (input_counter == 2) ? -0x18bd : (input_counter == 3) ? -0x1e9f : (input_counter == 4) ? -0x94a : (input_counter == 5) ? 0x144d : (input_counter == 6) ? 0x1fd9 : (input_counter == 7) ? 0x0f16 : (input_counter == 8) ? -0xf16 : (input_counter == 9) ? -0x1fd9 : (input_counter == 10) ? -0x144d : (input_counter == 11) ? 0x094a : (input_counter == 12) ? 0x1e9f : (input_counter == 13) ? 0x18bd : (input_counter == 14) ? -0x323 : (input_counter == 15) ? -0x1c39 : (input_counter == 16) ? -0x1c39 : (input_counter == 17) ? -0x323 : (input_counter == 18) ? 0x18bd : (input_counter == 19) ? 0x1e9f : (input_counter == 20) ? 0x094a : (input_counter == 21) ? -0x144d : (input_counter == 22) ? -0x1fd9 : (input_counter == 23) ? -0xf16 : (input_counter == 24) ? 0x0f16 : (input_counter == 25) ? 0x1fd9 : (input_counter == 26) ? 0x144d : (input_counter == 27) ? -0x94a : (input_counter == 28) ? -0x1e9f : (input_counter == 29) ? -0x18bd : (input_counter == 30) ? 0x0323 : 0x1c39;
11: coeff = (input_counter == 0) ? 0x1b73 : (input_counter == 1) ? -0x192 : (input_counter == 2) ? -0x1ced : (input_counter == 3) ? -0x19b4 : (input_counter == 4) ? 0x04b2 : (input_counter == 5) ? 0x1e21 : (input_counter == 6) ? 0x17b6 : (input_counter == 7) ? -0x7c6 : (input_counter == 8) ? -0x1f0a : (input_counter == 9) ? -0x157d : (input_counter == 10) ? 0x0ac8 : (input_counter == 11) ? 0x1fa7 : (input_counter == 12) ? 0x1310 : (input_counter == 13) ? -0xdaf : (input_counter == 14) ? -0x1ff6 : (input_counter == 15) ? -0x1074 : (input_counter == 16) ? 0x1074 : (input_counter == 17) ? 0x1ff6 : (input_counter == 18) ? 0x0daf : (input_counter == 19) ? -0x1310 : (input_counter == 20) ? -0x1fa7 : (input_counter == 21) ? -0xac8 : (input_counter == 22) ? 0x157d : (input_counter == 23) ? 0x1f0a : (input_counter == 24) ? 0x07c6 : (input_counter == 25) ? -0x17b6 : (input_counter == 26) ? -0x1e21 : (input_counter == 27) ? -0x4b2 : (input_counter == 28) ? 0x19b4 : (input_counter == 29) ? 0x1ced : (input_counter == 30) ? 0x0192 : -0x1b73;
12: coeff = (input_counter == 0) ? 0x1a9b : (input_counter == 1) ? -0x63e : (input_counter == 2) ? -0x1f63 : (input_counter == 3) ? -0x11c7 : (input_counter == 4) ? 0x11c7 : (input_counter == 5) ? 0x1f63 : (input_counter == 6) ? 0x063e : (input_counter == 7) ? -0x1a9b : (input_counter == 8) ? -0x1a9b : (input_counter == 9) ? 0x063e : (input_counter == 10) ? 0x1f63 : (input_counter == 11) ? 0x11c7 : (input_counter == 12) ? -0x11c7 : (input_counter == 13) ? -0x1f63 : (input_counter == 14) ? -0x63e : (input_counter == 15) ? 0x1a9b : (input_counter == 16) ? 0x1a9b : (input_counter == 17) ? -0x63e : (input_counter == 18) ? -0x1f63 : (input_counter == 19) ? -0x11c7 : (input_counter == 20) ? 0x11c7 : (input_counter == 21) ? 0x1f63 : (input_counter == 22) ? 0x063e : (input_counter == 23) ? -0x1a9b : (input_counter == 24) ? -0x1a9b : (input_counter == 25) ? 0x063e : (input_counter == 26) ? 0x1f63 : (input_counter == 27) ? 0x11c7 : (input_counter == 28) ? -0x11c7 : (input_counter == 29) ? -0x1f63 : (input_counter == 30) ? -0x63e : 0x1a9b;
13: coeff = (input_counter == 0) ? 0x19b4 : (input_counter == 1) ? -0xac8 : (input_counter == 2) ? -0x1ff6 : (input_counter == 3) ? -0x7c6 : (input_counter == 4) ? 0x1b73 : (input_counter == 5) ? 0x17b6 : (input_counter == 6) ? -0xdaf : (input_counter == 7) ? -0x1fa7 : (input_counter == 8) ? -0x4b2 : (input_counter == 9) ? 0x1ced : (input_counter == 10) ? 0x157d : (input_counter == 11) ? -0x1074 : (input_counter == 12) ? -0x1f0a : (input_counter == 13) ? -0x192 : (input_counter == 14) ? 0x1e21 : (input_counter == 15) ? 0x1310 : (input_counter == 16) ? -0x1310 : (input_counter == 17) ? -0x1e21 : (input_counter == 18) ? 0x0192 : (input_counter == 19) ? 0x1f0a : (input_counter == 20) ? 0x1074 : (input_counter == 21) ? -0x157d : (input_counter == 22) ? -0x1ced : (input_counter == 23) ? 0x04b2 : (input_counter == 24) ? 0x1fa7 : (input_counter == 25) ? 0x0daf : (input_counter == 26) ? -0x17b6 : (input_counter == 27) ? -0x1b73 : (input_counter == 28) ? 0x07c6 : (input_counter == 29) ? 0x1ff6 : (input_counter == 30) ? 0x0ac8 : -0x19b4;
14: coeff = (input_counter == 0) ? 0x18bd : (input_counter == 1) ? -0xf16 : (input_counter == 2) ? -0x1e9f : (input_counter == 3) ? 0x0323 : (input_counter == 4) ? 0x1fd9 : (input_counter == 5) ? 0x094a : (input_counter == 6) ? -0x1c39 : (input_counter == 7) ? -0x144d : (input_counter == 8) ? 0x144d : (input_counter == 9) ? 0x1c39 : (input_counter == 10) ? -0x94a : (input_counter == 11) ? -0x1fd9 : (input_counter == 12) ? -0x323 : (input_counter == 13) ? 0x1e9f : (input_counter == 14) ? 0x0f16 : (input_counter == 15) ? -0x18bd : (input_counter == 16) ? -0x18bd : (input_counter == 17) ? 0x0f16 : (input_counter == 18) ? 0x1e9f : (input_counter == 19) ? -0x323 : (input_counter == 20) ? -0x1fd9 : (input_counter == 21) ? -0x94a : (input_counter == 22) ? 0x1c39 : (input_counter == 23) ? 0x144d : (input_counter == 24) ? -0x144d : (input_counter == 25) ? -0x1c39 : (input_counter == 26) ? 0x094a : (input_counter == 27) ? 0x1fd9 : (input_counter == 28) ? 0x0323 : (input_counter == 29) ? -0x1e9f : (input_counter == 30) ? -0xf16 : 0x18bd;
15: coeff = (input_counter == 0) ? 0x17b6 : (input_counter == 1) ? -0x1310 : (input_counter == 2) ? -0x1b73 : (input_counter == 3) ? 0x0daf : (input_counter == 4) ? 0x1e21 : (input_counter == 5) ? -0x7c6 : (input_counter == 6) ? -0x1fa7 : (input_counter == 7) ? 0x0192 : (input_counter == 8) ? 0x1ff6 : (input_counter == 9) ? 0x04b2 : (input_counter == 10) ? -0x1f0a : (input_counter == 11) ? -0xac8 : (input_counter == 12) ? 0x1ced : (input_counter == 13) ? 0x1074 : (input_counter == 14) ? -0x19b4 : (input_counter == 15) ? -0x157d : (input_counter == 16) ? 0x157d : (input_counter == 17) ? 0x19b4 : (input_counter == 18) ? -0x1074 : (input_counter == 19) ? -0x1ced : (input_counter == 20) ? 0x0ac8 : (input_counter == 21) ? 0x1f0a : (input_counter == 22) ? -0x4b2 : (input_counter == 23) ? -0x1ff6 : (input_counter == 24) ? -0x192 : (input_counter == 25) ? 0x1fa7 : (input_counter == 26) ? 0x07c6 : (input_counter == 27) ? -0x1e21 : (input_counter == 28) ? -0xdaf : (input_counter == 29) ? 0x1b73 : (input_counter == 30) ? 0x1310 : -0x17b6;
16: coeff = (input_counter == 0) ? 0x16a1 : (input_counter == 1) ? -0x16a1 : (input_counter == 2) ? -0x16a1 : (input_counter == 3) ? 0x16a1 : (input_counter == 4) ? 0x16a1 : (input_counter == 5) ? -0x16a1 : (input_counter == 6) ? -0x16a1 : (input_counter == 7) ? 0x16a1 : (input_counter == 8) ? 0x16a1 : (input_counter == 9) ? -0x16a1 : (input_counter == 10) ? -0x16a1 : (input_counter == 11) ? 0x16a1 : (input_counter == 12) ? 0x16a1 : (input_counter == 13) ? -0x16a1 : (input_counter == 14) ? -0x16a1 : (input_counter == 15) ? 0x16a1 : (input_counter == 16) ? 0x16a1 : (input_counter == 17) ? -0x16a1 : (input_counter == 18) ? -0x16a1 : (input_counter == 19) ? 0x16a1 : (input_counter == 20) ? 0x16a1 : (input_counter == 21) ? -0x16a1 : (input_counter == 22) ? -0x16a1 : (input_counter == 23) ? 0x16a1 : (input_counter == 24) ? 0x16a1 : (input_counter == 25) ? -0x16a1 : (input_counter == 26) ? -0x16a1 : (input_counter == 27) ? 0x16a1 : (input_counter == 28) ? 0x16a1 : (input_counter == 29) ? -0x16a1 : (input_counter == 30) ? -0x16a1 : 0x16a1;
17: coeff = (input_counter == 0) ? 0x157d : (input_counter == 1) ? -0x19b4 : (input_counter == 2) ? -0x1074 : (input_counter == 3) ? 0x1ced : (input_counter == 4) ? 0x0ac8 : (input_counter == 5) ? -0x1f0a : (input_counter == 6) ? -0x4b2 : (input_counter == 7) ? 0x1ff6 : (input_counter == 8) ? -0x192 : (input_counter == 9) ? -0x1fa7 : (input_counter == 10) ? 0x07c6 : (input_counter == 11) ? 0x1e21 : (input_counter == 12) ? -0xdaf : (input_counter == 13) ? -0x1b73 : (input_counter == 14) ? 0x1310 : (input_counter == 15) ? 0x17b6 : (input_counter == 16) ? -0x17b6 : (input_counter == 17) ? -0x1310 : (input_counter == 18) ? 0x1b73 : (input_counter == 19) ? 0x0daf : (input_counter == 20) ? -0x1e21 : (input_counter == 21) ? -0x7c6 : (input_counter == 22) ? 0x1fa7 : (input_counter == 23) ? 0x0192 : (input_counter == 24) ? -0x1ff6 : (input_counter == 25) ? 0x04b2 : (input_counter == 26) ? 0x1f0a : (input_counter == 27) ? -0xac8 : (input_counter == 28) ? -0x1ced : (input_counter == 29) ? 0x1074 : (input_counter == 30) ? 0x19b4 : -0x157d;
18: coeff = (input_counter == 0) ? 0x144d : (input_counter == 1) ? -0x1c39 : (input_counter == 2) ? -0x94a : (input_counter == 3) ? 0x1fd9 : (input_counter == 4) ? -0x323 : (input_counter == 5) ? -0x1e9f : (input_counter == 6) ? 0x0f16 : (input_counter == 7) ? 0x18bd : (input_counter == 8) ? -0x18bd : (input_counter == 9) ? -0xf16 : (input_counter == 10) ? 0x1e9f : (input_counter == 11) ? 0x0323 : (input_counter == 12) ? -0x1fd9 : (input_counter == 13) ? 0x094a : (input_counter == 14) ? 0x1c39 : (input_counter == 15) ? -0x144d : (input_counter == 16) ? -0x144d : (input_counter == 17) ? 0x1c39 : (input_counter == 18) ? 0x094a : (input_counter == 19) ? -0x1fd9 : (input_counter == 20) ? 0x0323 : (input_counter == 21) ? 0x1e9f : (input_counter == 22) ? -0xf16 : (input_counter == 23) ? -0x18bd : (input_counter == 24) ? 0x18bd : (input_counter == 25) ? 0x0f16 : (input_counter == 26) ? -0x1e9f : (input_counter == 27) ? -0x323 : (input_counter == 28) ? 0x1fd9 : (input_counter == 29) ? -0x94a : (input_counter == 30) ? -0x1c39 : 0x144d;
19: coeff = (input_counter == 0) ? 0x1310 : (input_counter == 1) ? -0x1e21 : (input_counter == 2) ? -0x192 : (input_counter == 3) ? 0x1f0a : (input_counter == 4) ? -0x1074 : (input_counter == 5) ? -0x157d : (input_counter == 6) ? 0x1ced : (input_counter == 7) ? 0x04b2 : (input_counter == 8) ? -0x1fa7 : (input_counter == 9) ? 0x0daf : (input_counter == 10) ? 0x17b6 : (input_counter == 11) ? -0x1b73 : (input_counter == 12) ? -0x7c6 : (input_counter == 13) ? 0x1ff6 : (input_counter == 14) ? -0xac8 : (input_counter == 15) ? -0x19b4 : (input_counter == 16) ? 0x19b4 : (input_counter == 17) ? 0x0ac8 : (input_counter == 18) ? -0x1ff6 : (input_counter == 19) ? 0x07c6 : (input_counter == 20) ? 0x1b73 : (input_counter == 21) ? -0x17b6 : (input_counter == 22) ? -0xdaf : (input_counter == 23) ? 0x1fa7 : (input_counter == 24) ? -0x4b2 : (input_counter == 25) ? -0x1ced : (input_counter == 26) ? 0x157d : (input_counter == 27) ? 0x1074 : (input_counter == 28) ? -0x1f0a : (input_counter == 29) ? 0x0192 : (input_counter == 30) ? 0x1e21 : -0x1310;
20: coeff = (input_counter == 0) ? 0x11c7 : (input_counter == 1) ? -0x1f63 : (input_counter == 2) ? 0x063e : (input_counter == 3) ? 0x1a9b : (input_counter == 4) ? -0x1a9b : (input_counter == 5) ? -0x63e : (input_counter == 6) ? 0x1f63 : (input_counter == 7) ? -0x11c7 : (input_counter == 8) ? -0x11c7 : (input_counter == 9) ? 0x1f63 : (input_counter == 10) ? -0x63e : (input_counter == 11) ? -0x1a9b : (input_counter == 12) ? 0x1a9b : (input_counter == 13) ? 0x063e : (input_counter == 14) ? -0x1f63 : (input_counter == 15) ? 0x11c7 : (input_counter == 16) ? 0x11c7 : (input_counter == 17) ? -0x1f63 : (input_counter == 18) ? 0x063e : (input_counter == 19) ? 0x1a9b : (input_counter == 20) ? -0x1a9b : (input_counter == 21) ? -0x63e : (input_counter == 22) ? 0x1f63 : (input_counter == 23) ? -0x11c7 : (input_counter == 24) ? -0x11c7 : (input_counter == 25) ? 0x1f63 : (input_counter == 26) ? -0x63e : (input_counter == 27) ? -0x1a9b : (input_counter == 28) ? 0x1a9b : (input_counter == 29) ? 0x063e : (input_counter == 30) ? -0x1f63 : 0x11c7;
21: coeff = (input_counter == 0) ? 0x1074 : (input_counter == 1) ? -0x1ff6 : (input_counter == 2) ? 0x0daf : (input_counter == 3) ? 0x1310 : (input_counter == 4) ? -0x1fa7 : (input_counter == 5) ? 0x0ac8 : (input_counter == 6) ? 0x157d : (input_counter == 7) ? -0x1f0a : (input_counter == 8) ? 0x07c6 : (input_counter == 9) ? 0x17b6 : (input_counter == 10) ? -0x1e21 : (input_counter == 11) ? 0x04b2 : (input_counter == 12) ? 0x19b4 : (input_counter == 13) ? -0x1ced : (input_counter == 14) ? 0x0192 : (input_counter == 15) ? 0x1b73 : (input_counter == 16) ? -0x1b73 : (input_counter == 17) ? -0x192 : (input_counter == 18) ? 0x1ced : (input_counter == 19) ? -0x19b4 : (input_counter == 20) ? -0x4b2 : (input_counter == 21) ? 0x1e21 : (input_counter == 22) ? -0x17b6 : (input_counter == 23) ? -0x7c6 : (input_counter == 24) ? 0x1f0a : (input_counter == 25) ? -0x157d : (input_counter == 26) ? -0xac8 : (input_counter == 27) ? 0x1fa7 : (input_counter == 28) ? -0x1310 : (input_counter == 29) ? -0xdaf : (input_counter == 30) ? 0x1ff6 : -0x1074;
22: coeff = (input_counter == 0) ? 0x0f16 : (input_counter == 1) ? -0x1fd9 : (input_counter == 2) ? 0x144d : (input_counter == 3) ? 0x094a : (input_counter == 4) ? -0x1e9f : (input_counter == 5) ? 0x18bd : (input_counter == 6) ? 0x0323 : (input_counter == 7) ? -0x1c39 : (input_counter == 8) ? 0x1c39 : (input_counter == 9) ? -0x323 : (input_counter == 10) ? -0x18bd : (input_counter == 11) ? 0x1e9f : (input_counter == 12) ? -0x94a : (input_counter == 13) ? -0x144d : (input_counter == 14) ? 0x1fd9 : (input_counter == 15) ? -0xf16 : (input_counter == 16) ? -0xf16 : (input_counter == 17) ? 0x1fd9 : (input_counter == 18) ? -0x144d : (input_counter == 19) ? -0x94a : (input_counter == 20) ? 0x1e9f : (input_counter == 21) ? -0x18bd : (input_counter == 22) ? -0x323 : (input_counter == 23) ? 0x1c39 : (input_counter == 24) ? -0x1c39 : (input_counter == 25) ? 0x0323 : (input_counter == 26) ? 0x18bd : (input_counter == 27) ? -0x1e9f : (input_counter == 28) ? 0x094a : (input_counter == 29) ? 0x144d : (input_counter == 30) ? -0x1fd9 : 0x0f16;
23: coeff = (input_counter == 0) ? 0x0daf : (input_counter == 1) ? -0x1f0a : (input_counter == 2) ? 0x19b4 : (input_counter == 3) ? -0x192 : (input_counter == 4) ? -0x17b6 : (input_counter == 5) ? 0x1fa7 : (input_counter == 6) ? -0x1074 : (input_counter == 7) ? -0xac8 : (input_counter == 8) ? 0x1e21 : (input_counter == 9) ? -0x1b73 : (input_counter == 10) ? 0x04b2 : (input_counter == 11) ? 0x157d : (input_counter == 12) ? -0x1ff6 : (input_counter == 13) ? 0x1310 : (input_counter == 14) ? 0x07c6 : (input_counter == 15) ? -0x1ced : (input_counter == 16) ? 0x1ced : (input_counter == 17) ? -0x7c6 : (input_counter == 18) ? -0x1310 : (input_counter == 19) ? 0x1ff6 : (input_counter == 20) ? -0x157d : (input_counter == 21) ? -0x4b2 : (input_counter == 22) ? 0x1b73 : (input_counter == 23) ? -0x1e21 : (input_counter == 24) ? 0x0ac8 : (input_counter == 25) ? 0x1074 : (input_counter == 26) ? -0x1fa7 : (input_counter == 27) ? 0x17b6 : (input_counter == 28) ? 0x0192 : (input_counter == 29) ? -0x19b4 : (input_counter == 30) ? 0x1f0a : -0xdaf;
24: coeff = (input_counter == 0) ? 0x0c3f : (input_counter == 1) ? -0x1d90 : (input_counter == 2) ? 0x1d90 : (input_counter == 3) ? -0xc3f : (input_counter == 4) ? -0xc3f : (input_counter == 5) ? 0x1d90 : (input_counter == 6) ? -0x1d90 : (input_counter == 7) ? 0x0c3f : (input_counter == 8) ? 0x0c3f : (input_counter == 9) ? -0x1d90 : (input_counter == 10) ? 0x1d90 : (input_counter == 11) ? -0xc3f : (input_counter == 12) ? -0xc3f : (input_counter == 13) ? 0x1d90 : (input_counter == 14) ? -0x1d90 : (input_counter == 15) ? 0x0c3f : (input_counter == 16) ? 0x0c3f : (input_counter == 17) ? -0x1d90 : (input_counter == 18) ? 0x1d90 : (input_counter == 19) ? -0xc3f : (input_counter == 20) ? -0xc3f : (input_counter == 21) ? 0x1d90 : (input_counter == 22) ? -0x1d90 : (input_counter == 23) ? 0x0c3f : (input_counter == 24) ? 0x0c3f : (input_counter == 25) ? -0x1d90 : (input_counter == 26) ? 0x1d90 : (input_counter == 27) ? -0xc3f : (input_counter == 28) ? -0xc3f : (input_counter == 29) ? 0x1d90 : (input_counter == 30) ? -0x1d90 : 0x0c3f;
25: coeff = (input_counter == 0) ? 0x0ac8 : (input_counter == 1) ? -0x1b73 : (input_counter == 2) ? 0x1fa7 : (input_counter == 3) ? -0x157d : (input_counter == 4) ? 0x0192 : (input_counter == 5) ? 0x1310 : (input_counter == 6) ? -0x1f0a : (input_counter == 7) ? 0x1ced : (input_counter == 8) ? -0xdaf : (input_counter == 9) ? -0x7c6 : (input_counter == 10) ? 0x19b4 : (input_counter == 11) ? -0x1ff6 : (input_counter == 12) ? 0x17b6 : (input_counter == 13) ? -0x4b2 : (input_counter == 14) ? -0x1074 : (input_counter == 15) ? 0x1e21 : (input_counter == 16) ? -0x1e21 : (input_counter == 17) ? 0x1074 : (input_counter == 18) ? 0x04b2 : (input_counter == 19) ? -0x17b6 : (input_counter == 20) ? 0x1ff6 : (input_counter == 21) ? -0x19b4 : (input_counter == 22) ? 0x07c6 : (input_counter == 23) ? 0x0daf : (input_counter == 24) ? -0x1ced : (input_counter == 25) ? 0x1f0a : (input_counter == 26) ? -0x1310 : (input_counter == 27) ? -0x192 : (input_counter == 28) ? 0x157d : (input_counter == 29) ? -0x1fa7 : (input_counter == 30) ? 0x1b73 : -0xac8;
26: coeff = (input_counter == 0) ? 0x094a : (input_counter == 1) ? -0x18bd : (input_counter == 2) ? 0x1fd9 : (input_counter == 3) ? -0x1c39 : (input_counter == 4) ? 0x0f16 : (input_counter == 5) ? 0x0323 : (input_counter == 6) ? -0x144d : (input_counter == 7) ? 0x1e9f : (input_counter == 8) ? -0x1e9f : (input_counter == 9) ? 0x144d : (input_counter == 10) ? -0x323 : (input_counter == 11) ? -0xf16 : (input_counter == 12) ? 0x1c39 : (input_counter == 13) ? -0x1fd9 : (input_counter == 14) ? 0x18bd : (input_counter == 15) ? -0x94a : (input_counter == 16) ? -0x94a : (input_counter == 17) ? 0x18bd : (input_counter == 18) ? -0x1fd9 : (input_counter == 19) ? 0x1c39 : (input_counter == 20) ? -0xf16 : (input_counter == 21) ? -0x323 : (input_counter == 22) ? 0x144d : (input_counter == 23) ? -0x1e9f : (input_counter == 24) ? 0x1e9f : (input_counter == 25) ? -0x144d : (input_counter == 26) ? 0x0323 : (input_counter == 27) ? 0x0f16 : (input_counter == 28) ? -0x1c39 : (input_counter == 29) ? 0x1fd9 : (input_counter == 30) ? -0x18bd : 0x094a;
27: coeff = (input_counter == 0) ? 0x07c6 : (input_counter == 1) ? -0x157d : (input_counter == 2) ? 0x1e21 : (input_counter == 3) ? -0x1fa7 : (input_counter == 4) ? 0x19b4 : (input_counter == 5) ? -0xdaf : (input_counter == 6) ? -0x192 : (input_counter == 7) ? 0x1074 : (input_counter == 8) ? -0x1b73 : (input_counter == 9) ? 0x1ff6 : (input_counter == 10) ? -0x1ced : (input_counter == 11) ? 0x1310 : (input_counter == 12) ? -0x4b2 : (input_counter == 13) ? -0xac8 : (input_counter == 14) ? 0x17b6 : (input_counter == 15) ? -0x1f0a : (input_counter == 16) ? 0x1f0a : (input_counter == 17) ? -0x17b6 : (input_counter == 18) ? 0x0ac8 : (input_counter == 19) ? 0x04b2 : (input_counter == 20) ? -0x1310 : (input_counter == 21) ? 0x1ced : (input_counter == 22) ? -0x1ff6 : (input_counter == 23) ? 0x1b73 : (input_counter == 24) ? -0x1074 : (input_counter == 25) ? 0x0192 : (input_counter == 26) ? 0x0daf : (input_counter == 27) ? -0x19b4 : (input_counter == 28) ? 0x1fa7 : (input_counter == 29) ? -0x1e21 : (input_counter == 30) ? 0x157d : -0x7c6;
28: coeff = (input_counter == 0) ? 0x063e : (input_counter == 1) ? -0x11c7 : (input_counter == 2) ? 0x1a9b : (input_counter == 3) ? -0x1f63 : (input_counter == 4) ? 0x1f63 : (input_counter == 5) ? -0x1a9b : (input_counter == 6) ? 0x11c7 : (input_counter == 7) ? -0x63e : (input_counter == 8) ? -0x63e : (input_counter == 9) ? 0x11c7 : (input_counter == 10) ? -0x1a9b : (input_counter == 11) ? 0x1f63 : (input_counter == 12) ? -0x1f63 : (input_counter == 13) ? 0x1a9b : (input_counter == 14) ? -0x11c7 : (input_counter == 15) ? 0x063e : (input_counter == 16) ? 0x063e : (input_counter == 17) ? -0x11c7 : (input_counter == 18) ? 0x1a9b : (input_counter == 19) ? -0x1f63 : (input_counter == 20) ? 0x1f63 : (input_counter == 21) ? -0x1a9b : (input_counter == 22) ? 0x11c7 : (input_counter == 23) ? -0x63e : (input_counter == 24) ? -0x63e : (input_counter == 25) ? 0x11c7 : (input_counter == 26) ? -0x1a9b : (input_counter == 27) ? 0x1f63 : (input_counter == 28) ? -0x1f63 : (input_counter == 29) ? 0x1a9b : (input_counter == 30) ? -0x11c7 : 0x063e;
29: coeff = (input_counter == 0) ? 0x04b2 : (input_counter == 1) ? -0xdaf : (input_counter == 2) ? 0x157d : (input_counter == 3) ? -0x1b73 : (input_counter == 4) ? 0x1f0a : (input_counter == 5) ? -0x1ff6 : (input_counter == 6) ? 0x1e21 : (input_counter == 7) ? -0x19b4 : (input_counter == 8) ? 0x1310 : (input_counter == 9) ? -0xac8 : (input_counter == 10) ? 0x0192 : (input_counter == 11) ? 0x07c6 : (input_counter == 12) ? -0x1074 : (input_counter == 13) ? 0x17b6 : (input_counter == 14) ? -0x1ced : (input_counter == 15) ? 0x1fa7 : (input_counter == 16) ? -0x1fa7 : (input_counter == 17) ? 0x1ced : (input_counter == 18) ? -0x17b6 : (input_counter == 19) ? 0x1074 : (input_counter == 20) ? -0x7c6 : (input_counter == 21) ? -0x192 : (input_counter == 22) ? 0x0ac8 : (input_counter == 23) ? -0x1310 : (input_counter == 24) ? 0x19b4 : (input_counter == 25) ? -0x1e21 : (input_counter == 26) ? 0x1ff6 : (input_counter == 27) ? -0x1f0a : (input_counter == 28) ? 0x1b73 : (input_counter == 29) ? -0x157d : (input_counter == 30) ? 0x0daf : -0x4b2;
30: coeff = (input_counter == 0) ? 0x0323 : (input_counter == 1) ? -0x94a : (input_counter == 2) ? 0x0f16 : (input_counter == 3) ? -0x144d : (input_counter == 4) ? 0x18bd : (input_counter == 5) ? -0x1c39 : (input_counter == 6) ? 0x1e9f : (input_counter == 7) ? -0x1fd9 : (input_counter == 8) ? 0x1fd9 : (input_counter == 9) ? -0x1e9f : (input_counter == 10) ? 0x1c39 : (input_counter == 11) ? -0x18bd : (input_counter == 12) ? 0x144d : (input_counter == 13) ? -0xf16 : (input_counter == 14) ? 0x094a : (input_counter == 15) ? -0x323 : (input_counter == 16) ? -0x323 : (input_counter == 17) ? 0x094a : (input_counter == 18) ? -0xf16 : (input_counter == 19) ? 0x144d : (input_counter == 20) ? -0x18bd : (input_counter == 21) ? 0x1c39 : (input_counter == 22) ? -0x1e9f : (input_counter == 23) ? 0x1fd9 : (input_counter == 24) ? -0x1fd9 : (input_counter == 25) ? 0x1e9f : (input_counter == 26) ? -0x1c39 : (input_counter == 27) ? 0x18bd : (input_counter == 28) ? -0x144d : (input_counter == 29) ? 0x0f16 : (input_counter == 30) ? -0x94a : 0x0323;
31: coeff = (input_counter == 0) ? 0x0192 : (input_counter == 1) ? -0x4b2 : (input_counter == 2) ? 0x07c6 : (input_counter == 3) ? -0xac8 : (input_counter == 4) ? 0x0daf : (input_counter == 5) ? -0x1074 : (input_counter == 6) ? 0x1310 : (input_counter == 7) ? -0x157d : (input_counter == 8) ? 0x17b6 : (input_counter == 9) ? -0x19b4 : (input_counter == 10) ? 0x1b73 : (input_counter == 11) ? -0x1ced : (input_counter == 12) ? 0x1e21 : (input_counter == 13) ? -0x1f0a : (input_counter == 14) ? 0x1fa7 : (input_counter == 15) ? -0x1ff6 : (input_counter == 16) ? 0x1ff6 : (input_counter == 17) ? -0x1fa7 : (input_counter == 18) ? 0x1f0a : (input_counter == 19) ? -0x1e21 : (input_counter == 20) ? 0x1ced : (input_counter == 21) ? -0x1b73 : (input_counter == 22) ? 0x19b4 : (input_counter == 23) ? -0x17b6 : (input_counter == 24) ? 0x157d : (input_counter == 25) ? -0x1310 : (input_counter == 26) ? 0x1074 : (input_counter == 27) ? -0xdaf : (input_counter == 28) ? 0x0ac8 : (input_counter == 29) ? -0x7c6 : (input_counter == 30) ? 0x04b2 : -0x192;
      default: coeff = 16'h0000;
    endcase
  end

   always @(posedge clk) begin
    if (rst) begin
      input_counter <= 0;
      output_counter <= 0;
      accumulator <= 0;
      dct_out <= 0;
      dct_valid <= 0;
      state <= 0;
    end else begin
      case (state)
        0: begin
          if (data_valid) begin
            input_buffer[input_counter] <= data_in;
            input_counter <= input_counter + 1;
            if (input_counter == N - 1) begin
              input_counter <= 0;
              state <= 1;
            end
          end
        end

        1: begin
          coeff <= dct_coeff(output_counter, input_counter);
          mult <= input_buffer[input_counter] * coeff;
          accumulator <= accumulator + mult;
          input_counter <= input_counter + 1;

          if (input_counter == N - 1) begin
            dct_out <= accumulator >>> (Q_L + COEFF_WIDTH - Q_D);
            dct_valid <= 1;
            accumulator <= 0;
            output_counter <= output_counter + 1;
            input_counter <= 0;

            if (output_counter == N - 1) begin
              output_counter <= 0;
              state <= 0;
            end
          end
        end
      endcase
    end
  end

endmodule

endmodule
`ifndef MEL_FILTERBANK_V
`define MEL_FILTERBANK_V

module mel_filterbank #(
    parameter NUM_MEL_FILTERS = 40,
    parameter NUM_DFT_POINTS = 256,
    parameter COEF_WIDTH = 16,
    parameter ACCUMULATOR_WIDTH = 32
) (
    input wire clk,
    input wire rst_n,
    input wire [31:0] dft_out,
    input wire dft_valid,
    output reg [ACCUMULATOR_WIDTH-1:0] mel_fbank_out,
    output reg mel_fbank_valid
);

    // Mel-scale filter coefficients (stored in LUT)
    reg [COEF_WIDTH-1:0] mel_filter_coefs [0:NUM_MEL_FILTERS-1][0:NUM_DFT_POINTS-1];

    // Registers for accumulating filterbank energies
    reg [ACCUMULATOR_WIDTH-1:0] mel_accumulators [0:NUM_MEL_FILTERS-1];

    // Counters for iterating over mel-scale filters and DFT points
    reg [$clog2(NUM_MEL_FILTERS)-1:0] mel_filter_cnt;
    reg [$clog2(NUM_DFT_POINTS)-1:0] dft_point_cnt;

  // Initialize mel-scale filter coefficients (precomputed)
    initial begin
	mel_filter_coefs[0][0] = 16'h0000;
	mel_filter_coefs[0][1] = 16'h5A7F;
	mel_filter_coefs[0][2] = 16'h4E2B;
	mel_filter_coefs[0][3] = 16'h0000;
	mel_filter_coefs[0][4] = 16'h0000;
	mel_filter_coefs[0][5] = 16'h0000;
	mel_filter_coefs[0][6] = 16'h0000;
	mel_filter_coefs[0][7] = 16'h0000;
	mel_filter_coefs[0][8] = 16'h0000;
	mel_filter_coefs[0][9] = 16'h0000;
	mel_filter_coefs[0][10] = 16'h0000;
	mel_filter_coefs[0][11] = 16'h0000;
	mel_filter_coefs[0][12] = 16'h0000;
	mel_filter_coefs[0][13] = 16'h0000;
	mel_filter_coefs[0][14] = 16'h0000;
	mel_filter_coefs[0][15] = 16'h0000;
	mel_filter_coefs[0][16] = 16'h0000;
	mel_filter_coefs[0][17] = 16'h0000;
	mel_filter_coefs[0][18] = 16'h0000;
	mel_filter_coefs[0][19] = 16'h0000;
	mel_filter_coefs[0][20] = 16'h0000;
	mel_filter_coefs[0][21] = 16'h0000;
	mel_filter_coefs[0][22] = 16'h0000;
	mel_filter_coefs[0][23] = 16'h0000;
	mel_filter_coefs[0][24] = 16'h0000;
	mel_filter_coefs[0][25] = 16'h0000;
	mel_filter_coefs[0][26] = 16'h0000;
	mel_filter_coefs[0][27] = 16'h0000;
	mel_filter_coefs[0][28] = 16'h0000;
	mel_filter_coefs[0][29] = 16'h0000;
	mel_filter_coefs[0][30] = 16'h0000;
	mel_filter_coefs[0][31] = 16'h0000;
	mel_filter_coefs[0][32] = 16'h0000;
	mel_filter_coefs[0][33] = 16'h0000;
	mel_filter_coefs[0][34] = 16'h0000;
	mel_filter_coefs[0][35] = 16'h0000;
	mel_filter_coefs[0][36] = 16'h0000;
	mel_filter_coefs[0][37] = 16'h0000;
	mel_filter_coefs[0][38] = 16'h0000;
	mel_filter_coefs[0][39] = 16'h0000;
	mel_filter_coefs[0][40] = 16'h0000;
	mel_filter_coefs[0][41] = 16'h0000;
	mel_filter_coefs[0][42] = 16'h0000;
	mel_filter_coefs[0][43] = 16'h0000;
	mel_filter_coefs[0][44] = 16'h0000;
	mel_filter_coefs[0][45] = 16'h0000;
	mel_filter_coefs[0][46] = 16'h0000;
	mel_filter_coefs[0][47] = 16'h0000;
	mel_filter_coefs[0][48] = 16'h0000;
	mel_filter_coefs[0][49] = 16'h0000;
	mel_filter_coefs[0][50] = 16'h0000;
	mel_filter_coefs[0][51] = 16'h0000;
	mel_filter_coefs[0][52] = 16'h0000;
	mel_filter_coefs[0][53] = 16'h0000;
	mel_filter_coefs[0][54] = 16'h0000;
	mel_filter_coefs[0][55] = 16'h0000;
	mel_filter_coefs[0][56] = 16'h0000;
	mel_filter_coefs[0][57] = 16'h0000;
	mel_filter_coefs[0][58] = 16'h0000;
	mel_filter_coefs[0][59] = 16'h0000;
	mel_filter_coefs[0][60] = 16'h0000;
	mel_filter_coefs[0][61] = 16'h0000;
	mel_filter_coefs[0][62] = 16'h0000;
	mel_filter_coefs[0][63] = 16'h0000;
	mel_filter_coefs[0][64] = 16'h0000;
	mel_filter_coefs[0][65] = 16'h0000;
	mel_filter_coefs[0][66] = 16'h0000;
	mel_filter_coefs[0][67] = 16'h0000;
	mel_filter_coefs[0][68] = 16'h0000;
	mel_filter_coefs[0][69] = 16'h0000;
	mel_filter_coefs[0][70] = 16'h0000;
	mel_filter_coefs[0][71] = 16'h0000;
	mel_filter_coefs[0][72] = 16'h0000;
	mel_filter_coefs[0][73] = 16'h0000;
	mel_filter_coefs[0][74] = 16'h0000;
	mel_filter_coefs[0][75] = 16'h0000;
	mel_filter_coefs[0][76] = 16'h0000;
	mel_filter_coefs[0][77] = 16'h0000;
	mel_filter_coefs[0][78] = 16'h0000;
	mel_filter_coefs[0][79] = 16'h0000;
	mel_filter_coefs[0][80] = 16'h0000;
	mel_filter_coefs[0][81] = 16'h0000;
	mel_filter_coefs[0][82] = 16'h0000;
	mel_filter_coefs[0][83] = 16'h0000;
	mel_filter_coefs[0][84] = 16'h0000;
	mel_filter_coefs[0][85] = 16'h0000;
	mel_filter_coefs[0][86] = 16'h0000;
	mel_filter_coefs[0][87] = 16'h0000;
	mel_filter_coefs[0][88] = 16'h0000;
	mel_filter_coefs[0][89] = 16'h0000;
	mel_filter_coefs[0][90] = 16'h0000;
	mel_filter_coefs[0][91] = 16'h0000;
	mel_filter_coefs[0][92] = 16'h0000;
	mel_filter_coefs[0][93] = 16'h0000;
	mel_filter_coefs[0][94] = 16'h0000;
	mel_filter_coefs[0][95] = 16'h0000;
	mel_filter_coefs[0][96] = 16'h0000;
	mel_filter_coefs[0][97] = 16'h0000;
	mel_filter_coefs[0][98] = 16'h0000;
	mel_filter_coefs[0][99] = 16'h0000;
	mel_filter_coefs[0][100] = 16'h0000;
	mel_filter_coefs[0][101] = 16'h0000;
	mel_filter_coefs[0][102] = 16'h0000;
	mel_filter_coefs[0][103] = 16'h0000;
	mel_filter_coefs[0][104] = 16'h0000;
	mel_filter_coefs[0][105] = 16'h0000;
	mel_filter_coefs[0][106] = 16'h0000;
	mel_filter_coefs[0][107] = 16'h0000;
	mel_filter_coefs[0][108] = 16'h0000;
	mel_filter_coefs[0][109] = 16'h0000;
	mel_filter_coefs[0][110] = 16'h0000;
	mel_filter_coefs[0][111] = 16'h0000;
	mel_filter_coefs[0][112] = 16'h0000;
	mel_filter_coefs[0][113] = 16'h0000;
	mel_filter_coefs[0][114] = 16'h0000;
	mel_filter_coefs[0][115] = 16'h0000;
	mel_filter_coefs[0][116] = 16'h0000;
	mel_filter_coefs[0][117] = 16'h0000;
	mel_filter_coefs[0][118] = 16'h0000;
	mel_filter_coefs[0][119] = 16'h0000;
	mel_filter_coefs[0][120] = 16'h0000;
	mel_filter_coefs[0][121] = 16'h0000;
	mel_filter_coefs[0][122] = 16'h0000;
	mel_filter_coefs[0][123] = 16'h0000;
	mel_filter_coefs[0][124] = 16'h0000;
	mel_filter_coefs[0][125] = 16'h0000;
	mel_filter_coefs[0][126] = 16'h0000;
	mel_filter_coefs[0][127] = 16'h0000;
	mel_filter_coefs[0][128] = 16'h0000;
	mel_filter_coefs[0][129] = 16'h0000;
	mel_filter_coefs[0][130] = 16'h0000;
	mel_filter_coefs[0][131] = 16'h0000;
	mel_filter_coefs[0][132] = 16'h0000;
	mel_filter_coefs[0][133] = 16'h0000;
	mel_filter_coefs[0][134] = 16'h0000;
	mel_filter_coefs[0][135] = 16'h0000;
	mel_filter_coefs[0][136] = 16'h0000;
	mel_filter_coefs[0][137] = 16'h0000;
	mel_filter_coefs[0][138] = 16'h0000;
	mel_filter_coefs[0][139] = 16'h0000;
	mel_filter_coefs[0][140] = 16'h0000;
	mel_filter_coefs[0][141] = 16'h0000;
	mel_filter_coefs[0][142] = 16'h0000;
	mel_filter_coefs[0][143] = 16'h0000;
	mel_filter_coefs[0][144] = 16'h0000;
	mel_filter_coefs[0][145] = 16'h0000;
	mel_filter_coefs[0][146] = 16'h0000;
	mel_filter_coefs[0][147] = 16'h0000;
	mel_filter_coefs[0][148] = 16'h0000;
	mel_filter_coefs[0][149] = 16'h0000;
	mel_filter_coefs[0][150] = 16'h0000;
	mel_filter_coefs[0][151] = 16'h0000;
	mel_filter_coefs[0][152] = 16'h0000;
	mel_filter_coefs[0][153] = 16'h0000;
	mel_filter_coefs[0][154] = 16'h0000;
	mel_filter_coefs[0][155] = 16'h0000;
	mel_filter_coefs[0][156] = 16'h0000;
	mel_filter_coefs[0][157] = 16'h0000;
	mel_filter_coefs[0][158] = 16'h0000;
	mel_filter_coefs[0][159] = 16'h0000;
	mel_filter_coefs[0][160] = 16'h0000;
	mel_filter_coefs[0][161] = 16'h0000;
	mel_filter_coefs[0][162] = 16'h0000;
	mel_filter_coefs[0][163] = 16'h0000;
	mel_filter_coefs[0][164] = 16'h0000;
	mel_filter_coefs[0][165] = 16'h0000;
	mel_filter_coefs[0][166] = 16'h0000;
	mel_filter_coefs[0][167] = 16'h0000;
	mel_filter_coefs[0][168] = 16'h0000;
	mel_filter_coefs[0][169] = 16'h0000;
	mel_filter_coefs[0][170] = 16'h0000;
	mel_filter_coefs[0][171] = 16'h0000;
	mel_filter_coefs[0][172] = 16'h0000;
	mel_filter_coefs[0][173] = 16'h0000;
	mel_filter_coefs[0][174] = 16'h0000;
	mel_filter_coefs[0][175] = 16'h0000;
	mel_filter_coefs[0][176] = 16'h0000;
	mel_filter_coefs[0][177] = 16'h0000;
	mel_filter_coefs[0][178] = 16'h0000;
	mel_filter_coefs[0][179] = 16'h0000;
	mel_filter_coefs[0][180] = 16'h0000;
	mel_filter_coefs[0][181] = 16'h0000;
	mel_filter_coefs[0][182] = 16'h0000;
	mel_filter_coefs[0][183] = 16'h0000;
	mel_filter_coefs[0][184] = 16'h0000;
	mel_filter_coefs[0][185] = 16'h0000;
	mel_filter_coefs[0][186] = 16'h0000;
	mel_filter_coefs[0][187] = 16'h0000;
	mel_filter_coefs[0][188] = 16'h0000;
	mel_filter_coefs[0][189] = 16'h0000;
	mel_filter_coefs[0][190] = 16'h0000;
	mel_filter_coefs[0][191] = 16'h0000;
	mel_filter_coefs[0][192] = 16'h0000;
	mel_filter_coefs[0][193] = 16'h0000;
	mel_filter_coefs[0][194] = 16'h0000;
	mel_filter_coefs[0][195] = 16'h0000;
	mel_filter_coefs[0][196] = 16'h0000;
	mel_filter_coefs[0][197] = 16'h0000;
	mel_filter_coefs[0][198] = 16'h0000;
	mel_filter_coefs[0][199] = 16'h0000;
	mel_filter_coefs[0][200] = 16'h0000;
	mel_filter_coefs[0][201] = 16'h0000;
	mel_filter_coefs[0][202] = 16'h0000;
	mel_filter_coefs[0][203] = 16'h0000;
	mel_filter_coefs[0][204] = 16'h0000;
	mel_filter_coefs[0][205] = 16'h0000;
	mel_filter_coefs[0][206] = 16'h0000;
	mel_filter_coefs[0][207] = 16'h0000;
	mel_filter_coefs[0][208] = 16'h0000;
	mel_filter_coefs[0][209] = 16'h0000;
	mel_filter_coefs[0][210] = 16'h0000;
	mel_filter_coefs[0][211] = 16'h0000;
	mel_filter_coefs[0][212] = 16'h0000;
	mel_filter_coefs[0][213] = 16'h0000;
	mel_filter_coefs[0][214] = 16'h0000;
	mel_filter_coefs[0][215] = 16'h0000;
	mel_filter_coefs[0][216] = 16'h0000;
	mel_filter_coefs[0][217] = 16'h0000;
	mel_filter_coefs[0][218] = 16'h0000;
	mel_filter_coefs[0][219] = 16'h0000;
	mel_filter_coefs[0][220] = 16'h0000;
	mel_filter_coefs[0][221] = 16'h0000;
	mel_filter_coefs[0][222] = 16'h0000;
	mel_filter_coefs[0][223] = 16'h0000;
	mel_filter_coefs[0][224] = 16'h0000;
	mel_filter_coefs[0][225] = 16'h0000;
	mel_filter_coefs[0][226] = 16'h0000;
	mel_filter_coefs[0][227] = 16'h0000;
	mel_filter_coefs[0][228] = 16'h0000;
	mel_filter_coefs[0][229] = 16'h0000;
	mel_filter_coefs[0][230] = 16'h0000;
	mel_filter_coefs[0][231] = 16'h0000;
	mel_filter_coefs[0][232] = 16'h0000;
	mel_filter_coefs[0][233] = 16'h0000;
	mel_filter_coefs[0][234] = 16'h0000;
	mel_filter_coefs[0][235] = 16'h0000;
	mel_filter_coefs[0][236] = 16'h0000;
	mel_filter_coefs[0][237] = 16'h0000;
	mel_filter_coefs[0][238] = 16'h0000;
	mel_filter_coefs[0][239] = 16'h0000;
	mel_filter_coefs[0][240] = 16'h0000;
	mel_filter_coefs[0][241] = 16'h0000;
	mel_filter_coefs[0][242] = 16'h0000;
	mel_filter_coefs[0][243] = 16'h0000;
	mel_filter_coefs[0][244] = 16'h0000;
	mel_filter_coefs[0][245] = 16'h0000;
	mel_filter_coefs[0][246] = 16'h0000;
	mel_filter_coefs[0][247] = 16'h0000;
	mel_filter_coefs[0][248] = 16'h0000;
	mel_filter_coefs[0][249] = 16'h0000;
	mel_filter_coefs[0][250] = 16'h0000;
	mel_filter_coefs[0][251] = 16'h0000;
	mel_filter_coefs[0][252] = 16'h0000;
	mel_filter_coefs[0][253] = 16'h0000;
	mel_filter_coefs[0][254] = 16'h0000;
	mel_filter_coefs[0][255] = 16'h0000;
	mel_filter_coefs[1][0] = 16'h0000;
	mel_filter_coefs[1][1] = 16'h0000;
	mel_filter_coefs[1][2] = 16'h31D5;
	mel_filter_coefs[1][3] = 16'h797A;
	mel_filter_coefs[1][4] = 16'h2973;
	mel_filter_coefs[1][5] = 16'h0000;
	mel_filter_coefs[1][6] = 16'h0000;
	mel_filter_coefs[1][7] = 16'h0000;
	mel_filter_coefs[1][8] = 16'h0000;
	mel_filter_coefs[1][9] = 16'h0000;
	mel_filter_coefs[1][10] = 16'h0000;
	mel_filter_coefs[1][11] = 16'h0000;
	mel_filter_coefs[1][12] = 16'h0000;
	mel_filter_coefs[1][13] = 16'h0000;
	mel_filter_coefs[1][14] = 16'h0000;
	mel_filter_coefs[1][15] = 16'h0000;
	mel_filter_coefs[1][16] = 16'h0000;
	mel_filter_coefs[1][17] = 16'h0000;
	mel_filter_coefs[1][18] = 16'h0000;
	mel_filter_coefs[1][19] = 16'h0000;
	mel_filter_coefs[1][20] = 16'h0000;
	mel_filter_coefs[1][21] = 16'h0000;
	mel_filter_coefs[1][22] = 16'h0000;
	mel_filter_coefs[1][23] = 16'h0000;
	mel_filter_coefs[1][24] = 16'h0000;
	mel_filter_coefs[1][25] = 16'h0000;
	mel_filter_coefs[1][26] = 16'h0000;
	mel_filter_coefs[1][27] = 16'h0000;
	mel_filter_coefs[1][28] = 16'h0000;
	mel_filter_coefs[1][29] = 16'h0000;
	mel_filter_coefs[1][30] = 16'h0000;
	mel_filter_coefs[1][31] = 16'h0000;
	mel_filter_coefs[1][32] = 16'h0000;
	mel_filter_coefs[1][33] = 16'h0000;
	mel_filter_coefs[1][34] = 16'h0000;
	mel_filter_coefs[1][35] = 16'h0000;
	mel_filter_coefs[1][36] = 16'h0000;
	mel_filter_coefs[1][37] = 16'h0000;
	mel_filter_coefs[1][38] = 16'h0000;
	mel_filter_coefs[1][39] = 16'h0000;
	mel_filter_coefs[1][40] = 16'h0000;
	mel_filter_coefs[1][41] = 16'h0000;
	mel_filter_coefs[1][42] = 16'h0000;
	mel_filter_coefs[1][43] = 16'h0000;
	mel_filter_coefs[1][44] = 16'h0000;
	mel_filter_coefs[1][45] = 16'h0000;
	mel_filter_coefs[1][46] = 16'h0000;
	mel_filter_coefs[1][47] = 16'h0000;
	mel_filter_coefs[1][48] = 16'h0000;
	mel_filter_coefs[1][49] = 16'h0000;
	mel_filter_coefs[1][50] = 16'h0000;
	mel_filter_coefs[1][51] = 16'h0000;
	mel_filter_coefs[1][52] = 16'h0000;
	mel_filter_coefs[1][53] = 16'h0000;
	mel_filter_coefs[1][54] = 16'h0000;
	mel_filter_coefs[1][55] = 16'h0000;
	mel_filter_coefs[1][56] = 16'h0000;
	mel_filter_coefs[1][57] = 16'h0000;
	mel_filter_coefs[1][58] = 16'h0000;
	mel_filter_coefs[1][59] = 16'h0000;
	mel_filter_coefs[1][60] = 16'h0000;
	mel_filter_coefs[1][61] = 16'h0000;
	mel_filter_coefs[1][62] = 16'h0000;
	mel_filter_coefs[1][63] = 16'h0000;
	mel_filter_coefs[1][64] = 16'h0000;
	mel_filter_coefs[1][65] = 16'h0000;
	mel_filter_coefs[1][66] = 16'h0000;
	mel_filter_coefs[1][67] = 16'h0000;
	mel_filter_coefs[1][68] = 16'h0000;
	mel_filter_coefs[1][69] = 16'h0000;
	mel_filter_coefs[1][70] = 16'h0000;
	mel_filter_coefs[1][71] = 16'h0000;
	mel_filter_coefs[1][72] = 16'h0000;
	mel_filter_coefs[1][73] = 16'h0000;
	mel_filter_coefs[1][74] = 16'h0000;
	mel_filter_coefs[1][75] = 16'h0000;
	mel_filter_coefs[1][76] = 16'h0000;
	mel_filter_coefs[1][77] = 16'h0000;
	mel_filter_coefs[1][78] = 16'h0000;
	mel_filter_coefs[1][79] = 16'h0000;
	mel_filter_coefs[1][80] = 16'h0000;
	mel_filter_coefs[1][81] = 16'h0000;
	mel_filter_coefs[1][82] = 16'h0000;
	mel_filter_coefs[1][83] = 16'h0000;
	mel_filter_coefs[1][84] = 16'h0000;
	mel_filter_coefs[1][85] = 16'h0000;
	mel_filter_coefs[1][86] = 16'h0000;
	mel_filter_coefs[1][87] = 16'h0000;
	mel_filter_coefs[1][88] = 16'h0000;
	mel_filter_coefs[1][89] = 16'h0000;
	mel_filter_coefs[1][90] = 16'h0000;
	mel_filter_coefs[1][91] = 16'h0000;
	mel_filter_coefs[1][92] = 16'h0000;
	mel_filter_coefs[1][93] = 16'h0000;
	mel_filter_coefs[1][94] = 16'h0000;
	mel_filter_coefs[1][95] = 16'h0000;
	mel_filter_coefs[1][96] = 16'h0000;
	mel_filter_coefs[1][97] = 16'h0000;
	mel_filter_coefs[1][98] = 16'h0000;
	mel_filter_coefs[1][99] = 16'h0000;
	mel_filter_coefs[1][100] = 16'h0000;
	mel_filter_coefs[1][101] = 16'h0000;
	mel_filter_coefs[1][102] = 16'h0000;
	mel_filter_coefs[1][103] = 16'h0000;
	mel_filter_coefs[1][104] = 16'h0000;
	mel_filter_coefs[1][105] = 16'h0000;
	mel_filter_coefs[1][106] = 16'h0000;
	mel_filter_coefs[1][107] = 16'h0000;
	mel_filter_coefs[1][108] = 16'h0000;
	mel_filter_coefs[1][109] = 16'h0000;
	mel_filter_coefs[1][110] = 16'h0000;
	mel_filter_coefs[1][111] = 16'h0000;
	mel_filter_coefs[1][112] = 16'h0000;
	mel_filter_coefs[1][113] = 16'h0000;
	mel_filter_coefs[1][114] = 16'h0000;
	mel_filter_coefs[1][115] = 16'h0000;
	mel_filter_coefs[1][116] = 16'h0000;
	mel_filter_coefs[1][117] = 16'h0000;
	mel_filter_coefs[1][118] = 16'h0000;
	mel_filter_coefs[1][119] = 16'h0000;
	mel_filter_coefs[1][120] = 16'h0000;
	mel_filter_coefs[1][121] = 16'h0000;
	mel_filter_coefs[1][122] = 16'h0000;
	mel_filter_coefs[1][123] = 16'h0000;
	mel_filter_coefs[1][124] = 16'h0000;
	mel_filter_coefs[1][125] = 16'h0000;
	mel_filter_coefs[1][126] = 16'h0000;
	mel_filter_coefs[1][127] = 16'h0000;
	mel_filter_coefs[1][128] = 16'h0000;
	mel_filter_coefs[1][129] = 16'h0000;
	mel_filter_coefs[1][130] = 16'h0000;
	mel_filter_coefs[1][131] = 16'h0000;
	mel_filter_coefs[1][132] = 16'h0000;
	mel_filter_coefs[1][133] = 16'h0000;
	mel_filter_coefs[1][134] = 16'h0000;
	mel_filter_coefs[1][135] = 16'h0000;
	mel_filter_coefs[1][136] = 16'h0000;
	mel_filter_coefs[1][137] = 16'h0000;
	mel_filter_coefs[1][138] = 16'h0000;
	mel_filter_coefs[1][139] = 16'h0000;
	mel_filter_coefs[1][140] = 16'h0000;
	mel_filter_coefs[1][141] = 16'h0000;
	mel_filter_coefs[1][142] = 16'h0000;
	mel_filter_coefs[1][143] = 16'h0000;
	mel_filter_coefs[1][144] = 16'h0000;
	mel_filter_coefs[1][145] = 16'h0000;
	mel_filter_coefs[1][146] = 16'h0000;
	mel_filter_coefs[1][147] = 16'h0000;
	mel_filter_coefs[1][148] = 16'h0000;
	mel_filter_coefs[1][149] = 16'h0000;
	mel_filter_coefs[1][150] = 16'h0000;
	mel_filter_coefs[1][151] = 16'h0000;
	mel_filter_coefs[1][152] = 16'h0000;
	mel_filter_coefs[1][153] = 16'h0000;
	mel_filter_coefs[1][154] = 16'h0000;
	mel_filter_coefs[1][155] = 16'h0000;
	mel_filter_coefs[1][156] = 16'h0000;
	mel_filter_coefs[1][157] = 16'h0000;
	mel_filter_coefs[1][158] = 16'h0000;
	mel_filter_coefs[1][159] = 16'h0000;
	mel_filter_coefs[1][160] = 16'h0000;
	mel_filter_coefs[1][161] = 16'h0000;
	mel_filter_coefs[1][162] = 16'h0000;
	mel_filter_coefs[1][163] = 16'h0000;
	mel_filter_coefs[1][164] = 16'h0000;
	mel_filter_coefs[1][165] = 16'h0000;
	mel_filter_coefs[1][166] = 16'h0000;
	mel_filter_coefs[1][167] = 16'h0000;
	mel_filter_coefs[1][168] = 16'h0000;
	mel_filter_coefs[1][169] = 16'h0000;
	mel_filter_coefs[1][170] = 16'h0000;
	mel_filter_coefs[1][171] = 16'h0000;
	mel_filter_coefs[1][172] = 16'h0000;
	mel_filter_coefs[1][173] = 16'h0000;
	mel_filter_coefs[1][174] = 16'h0000;
	mel_filter_coefs[1][175] = 16'h0000;
	mel_filter_coefs[1][176] = 16'h0000;
	mel_filter_coefs[1][177] = 16'h0000;
	mel_filter_coefs[1][178] = 16'h0000;
	mel_filter_coefs[1][179] = 16'h0000;
	mel_filter_coefs[1][180] = 16'h0000;
	mel_filter_coefs[1][181] = 16'h0000;
	mel_filter_coefs[1][182] = 16'h0000;
	mel_filter_coefs[1][183] = 16'h0000;
	mel_filter_coefs[1][184] = 16'h0000;
	mel_filter_coefs[1][185] = 16'h0000;
	mel_filter_coefs[1][186] = 16'h0000;
	mel_filter_coefs[1][187] = 16'h0000;
	mel_filter_coefs[1][188] = 16'h0000;
	mel_filter_coefs[1][189] = 16'h0000;
	mel_filter_coefs[1][190] = 16'h0000;
	mel_filter_coefs[1][191] = 16'h0000;
	mel_filter_coefs[1][192] = 16'h0000;
	mel_filter_coefs[1][193] = 16'h0000;
	mel_filter_coefs[1][194] = 16'h0000;
	mel_filter_coefs[1][195] = 16'h0000;
	mel_filter_coefs[1][196] = 16'h0000;
	mel_filter_coefs[1][197] = 16'h0000;
	mel_filter_coefs[1][198] = 16'h0000;
	mel_filter_coefs[1][199] = 16'h0000;
	mel_filter_coefs[1][200] = 16'h0000;
	mel_filter_coefs[1][201] = 16'h0000;
	mel_filter_coefs[1][202] = 16'h0000;
	mel_filter_coefs[1][203] = 16'h0000;
	mel_filter_coefs[1][204] = 16'h0000;
	mel_filter_coefs[1][205] = 16'h0000;
	mel_filter_coefs[1][206] = 16'h0000;
	mel_filter_coefs[1][207] = 16'h0000;
	mel_filter_coefs[1][208] = 16'h0000;
	mel_filter_coefs[1][209] = 16'h0000;
	mel_filter_coefs[1][210] = 16'h0000;
	mel_filter_coefs[1][211] = 16'h0000;
	mel_filter_coefs[1][212] = 16'h0000;
	mel_filter_coefs[1][213] = 16'h0000;
	mel_filter_coefs[1][214] = 16'h0000;
	mel_filter_coefs[1][215] = 16'h0000;
	mel_filter_coefs[1][216] = 16'h0000;
	mel_filter_coefs[1][217] = 16'h0000;
	mel_filter_coefs[1][218] = 16'h0000;
	mel_filter_coefs[1][219] = 16'h0000;
	mel_filter_coefs[1][220] = 16'h0000;
	mel_filter_coefs[1][221] = 16'h0000;
	mel_filter_coefs[1][222] = 16'h0000;
	mel_filter_coefs[1][223] = 16'h0000;
	mel_filter_coefs[1][224] = 16'h0000;
	mel_filter_coefs[1][225] = 16'h0000;
	mel_filter_coefs[1][226] = 16'h0000;
	mel_filter_coefs[1][227] = 16'h0000;
	mel_filter_coefs[1][228] = 16'h0000;
	mel_filter_coefs[1][229] = 16'h0000;
	mel_filter_coefs[1][230] = 16'h0000;
	mel_filter_coefs[1][231] = 16'h0000;
	mel_filter_coefs[1][232] = 16'h0000;
	mel_filter_coefs[1][233] = 16'h0000;
	mel_filter_coefs[1][234] = 16'h0000;
	mel_filter_coefs[1][235] = 16'h0000;
	mel_filter_coefs[1][236] = 16'h0000;
	mel_filter_coefs[1][237] = 16'h0000;
	mel_filter_coefs[1][238] = 16'h0000;
	mel_filter_coefs[1][239] = 16'h0000;
	mel_filter_coefs[1][240] = 16'h0000;
	mel_filter_coefs[1][241] = 16'h0000;
	mel_filter_coefs[1][242] = 16'h0000;
	mel_filter_coefs[1][243] = 16'h0000;
	mel_filter_coefs[1][244] = 16'h0000;
	mel_filter_coefs[1][245] = 16'h0000;
	mel_filter_coefs[1][246] = 16'h0000;
	mel_filter_coefs[1][247] = 16'h0000;
	mel_filter_coefs[1][248] = 16'h0000;
	mel_filter_coefs[1][249] = 16'h0000;
	mel_filter_coefs[1][250] = 16'h0000;
	mel_filter_coefs[1][251] = 16'h0000;
	mel_filter_coefs[1][252] = 16'h0000;
	mel_filter_coefs[1][253] = 16'h0000;
	mel_filter_coefs[1][254] = 16'h0000;
	mel_filter_coefs[1][255] = 16'h0000;
	mel_filter_coefs[2][0] = 16'h0000;
	mel_filter_coefs[2][1] = 16'h0000;
	mel_filter_coefs[2][2] = 16'h0000;
	mel_filter_coefs[2][3] = 16'h0686;
	mel_filter_coefs[2][4] = 16'h568D;
	mel_filter_coefs[2][5] = 16'h5BB9;
	mel_filter_coefs[2][6] = 16'h1077;
	mel_filter_coefs[2][7] = 16'h0000;
	mel_filter_coefs[2][8] = 16'h0000;
	mel_filter_coefs[2][9] = 16'h0000;
	mel_filter_coefs[2][10] = 16'h0000;
	mel_filter_coefs[2][11] = 16'h0000;
	mel_filter_coefs[2][12] = 16'h0000;
	mel_filter_coefs[2][13] = 16'h0000;
	mel_filter_coefs[2][14] = 16'h0000;
	mel_filter_coefs[2][15] = 16'h0000;
	mel_filter_coefs[2][16] = 16'h0000;
	mel_filter_coefs[2][17] = 16'h0000;
	mel_filter_coefs[2][18] = 16'h0000;
	mel_filter_coefs[2][19] = 16'h0000;
	mel_filter_coefs[2][20] = 16'h0000;
	mel_filter_coefs[2][21] = 16'h0000;
	mel_filter_coefs[2][22] = 16'h0000;
	mel_filter_coefs[2][23] = 16'h0000;
	mel_filter_coefs[2][24] = 16'h0000;
	mel_filter_coefs[2][25] = 16'h0000;
	mel_filter_coefs[2][26] = 16'h0000;
	mel_filter_coefs[2][27] = 16'h0000;
	mel_filter_coefs[2][28] = 16'h0000;
	mel_filter_coefs[2][29] = 16'h0000;
	mel_filter_coefs[2][30] = 16'h0000;
	mel_filter_coefs[2][31] = 16'h0000;
	mel_filter_coefs[2][32] = 16'h0000;
	mel_filter_coefs[2][33] = 16'h0000;
	mel_filter_coefs[2][34] = 16'h0000;
	mel_filter_coefs[2][35] = 16'h0000;
	mel_filter_coefs[2][36] = 16'h0000;
	mel_filter_coefs[2][37] = 16'h0000;
	mel_filter_coefs[2][38] = 16'h0000;
	mel_filter_coefs[2][39] = 16'h0000;
	mel_filter_coefs[2][40] = 16'h0000;
	mel_filter_coefs[2][41] = 16'h0000;
	mel_filter_coefs[2][42] = 16'h0000;
	mel_filter_coefs[2][43] = 16'h0000;
	mel_filter_coefs[2][44] = 16'h0000;
	mel_filter_coefs[2][45] = 16'h0000;
	mel_filter_coefs[2][46] = 16'h0000;
	mel_filter_coefs[2][47] = 16'h0000;
	mel_filter_coefs[2][48] = 16'h0000;
	mel_filter_coefs[2][49] = 16'h0000;
	mel_filter_coefs[2][50] = 16'h0000;
	mel_filter_coefs[2][51] = 16'h0000;
	mel_filter_coefs[2][52] = 16'h0000;
	mel_filter_coefs[2][53] = 16'h0000;
	mel_filter_coefs[2][54] = 16'h0000;
	mel_filter_coefs[2][55] = 16'h0000;
	mel_filter_coefs[2][56] = 16'h0000;
	mel_filter_coefs[2][57] = 16'h0000;
	mel_filter_coefs[2][58] = 16'h0000;
	mel_filter_coefs[2][59] = 16'h0000;
	mel_filter_coefs[2][60] = 16'h0000;
	mel_filter_coefs[2][61] = 16'h0000;
	mel_filter_coefs[2][62] = 16'h0000;
	mel_filter_coefs[2][63] = 16'h0000;
	mel_filter_coefs[2][64] = 16'h0000;
	mel_filter_coefs[2][65] = 16'h0000;
	mel_filter_coefs[2][66] = 16'h0000;
	mel_filter_coefs[2][67] = 16'h0000;
	mel_filter_coefs[2][68] = 16'h0000;
	mel_filter_coefs[2][69] = 16'h0000;
	mel_filter_coefs[2][70] = 16'h0000;
	mel_filter_coefs[2][71] = 16'h0000;
	mel_filter_coefs[2][72] = 16'h0000;
	mel_filter_coefs[2][73] = 16'h0000;
	mel_filter_coefs[2][74] = 16'h0000;
	mel_filter_coefs[2][75] = 16'h0000;
	mel_filter_coefs[2][76] = 16'h0000;
	mel_filter_coefs[2][77] = 16'h0000;
	mel_filter_coefs[2][78] = 16'h0000;
	mel_filter_coefs[2][79] = 16'h0000;
	mel_filter_coefs[2][80] = 16'h0000;
	mel_filter_coefs[2][81] = 16'h0000;
	mel_filter_coefs[2][82] = 16'h0000;
	mel_filter_coefs[2][83] = 16'h0000;
	mel_filter_coefs[2][84] = 16'h0000;
	mel_filter_coefs[2][85] = 16'h0000;
	mel_filter_coefs[2][86] = 16'h0000;
	mel_filter_coefs[2][87] = 16'h0000;
	mel_filter_coefs[2][88] = 16'h0000;
	mel_filter_coefs[2][89] = 16'h0000;
	mel_filter_coefs[2][90] = 16'h0000;
	mel_filter_coefs[2][91] = 16'h0000;
	mel_filter_coefs[2][92] = 16'h0000;
	mel_filter_coefs[2][93] = 16'h0000;
	mel_filter_coefs[2][94] = 16'h0000;
	mel_filter_coefs[2][95] = 16'h0000;
	mel_filter_coefs[2][96] = 16'h0000;
	mel_filter_coefs[2][97] = 16'h0000;
	mel_filter_coefs[2][98] = 16'h0000;
	mel_filter_coefs[2][99] = 16'h0000;
	mel_filter_coefs[2][100] = 16'h0000;
	mel_filter_coefs[2][101] = 16'h0000;
	mel_filter_coefs[2][102] = 16'h0000;
	mel_filter_coefs[2][103] = 16'h0000;
	mel_filter_coefs[2][104] = 16'h0000;
	mel_filter_coefs[2][105] = 16'h0000;
	mel_filter_coefs[2][106] = 16'h0000;
	mel_filter_coefs[2][107] = 16'h0000;
	mel_filter_coefs[2][108] = 16'h0000;
	mel_filter_coefs[2][109] = 16'h0000;
	mel_filter_coefs[2][110] = 16'h0000;
	mel_filter_coefs[2][111] = 16'h0000;
	mel_filter_coefs[2][112] = 16'h0000;
	mel_filter_coefs[2][113] = 16'h0000;
	mel_filter_coefs[2][114] = 16'h0000;
	mel_filter_coefs[2][115] = 16'h0000;
	mel_filter_coefs[2][116] = 16'h0000;
	mel_filter_coefs[2][117] = 16'h0000;
	mel_filter_coefs[2][118] = 16'h0000;
	mel_filter_coefs[2][119] = 16'h0000;
	mel_filter_coefs[2][120] = 16'h0000;
	mel_filter_coefs[2][121] = 16'h0000;
	mel_filter_coefs[2][122] = 16'h0000;
	mel_filter_coefs[2][123] = 16'h0000;
	mel_filter_coefs[2][124] = 16'h0000;
	mel_filter_coefs[2][125] = 16'h0000;
	mel_filter_coefs[2][126] = 16'h0000;
	mel_filter_coefs[2][127] = 16'h0000;
	mel_filter_coefs[2][128] = 16'h0000;
	mel_filter_coefs[2][129] = 16'h0000;
	mel_filter_coefs[2][130] = 16'h0000;
	mel_filter_coefs[2][131] = 16'h0000;
	mel_filter_coefs[2][132] = 16'h0000;
	mel_filter_coefs[2][133] = 16'h0000;
	mel_filter_coefs[2][134] = 16'h0000;
	mel_filter_coefs[2][135] = 16'h0000;
	mel_filter_coefs[2][136] = 16'h0000;
	mel_filter_coefs[2][137] = 16'h0000;
	mel_filter_coefs[2][138] = 16'h0000;
	mel_filter_coefs[2][139] = 16'h0000;
	mel_filter_coefs[2][140] = 16'h0000;
	mel_filter_coefs[2][141] = 16'h0000;
	mel_filter_coefs[2][142] = 16'h0000;
	mel_filter_coefs[2][143] = 16'h0000;
	mel_filter_coefs[2][144] = 16'h0000;
	mel_filter_coefs[2][145] = 16'h0000;
	mel_filter_coefs[2][146] = 16'h0000;
	mel_filter_coefs[2][147] = 16'h0000;
	mel_filter_coefs[2][148] = 16'h0000;
	mel_filter_coefs[2][149] = 16'h0000;
	mel_filter_coefs[2][150] = 16'h0000;
	mel_filter_coefs[2][151] = 16'h0000;
	mel_filter_coefs[2][152] = 16'h0000;
	mel_filter_coefs[2][153] = 16'h0000;
	mel_filter_coefs[2][154] = 16'h0000;
	mel_filter_coefs[2][155] = 16'h0000;
	mel_filter_coefs[2][156] = 16'h0000;
	mel_filter_coefs[2][157] = 16'h0000;
	mel_filter_coefs[2][158] = 16'h0000;
	mel_filter_coefs[2][159] = 16'h0000;
	mel_filter_coefs[2][160] = 16'h0000;
	mel_filter_coefs[2][161] = 16'h0000;
	mel_filter_coefs[2][162] = 16'h0000;
	mel_filter_coefs[2][163] = 16'h0000;
	mel_filter_coefs[2][164] = 16'h0000;
	mel_filter_coefs[2][165] = 16'h0000;
	mel_filter_coefs[2][166] = 16'h0000;
	mel_filter_coefs[2][167] = 16'h0000;
	mel_filter_coefs[2][168] = 16'h0000;
	mel_filter_coefs[2][169] = 16'h0000;
	mel_filter_coefs[2][170] = 16'h0000;
	mel_filter_coefs[2][171] = 16'h0000;
	mel_filter_coefs[2][172] = 16'h0000;
	mel_filter_coefs[2][173] = 16'h0000;
	mel_filter_coefs[2][174] = 16'h0000;
	mel_filter_coefs[2][175] = 16'h0000;
	mel_filter_coefs[2][176] = 16'h0000;
	mel_filter_coefs[2][177] = 16'h0000;
	mel_filter_coefs[2][178] = 16'h0000;
	mel_filter_coefs[2][179] = 16'h0000;
	mel_filter_coefs[2][180] = 16'h0000;
	mel_filter_coefs[2][181] = 16'h0000;
	mel_filter_coefs[2][182] = 16'h0000;
	mel_filter_coefs[2][183] = 16'h0000;
	mel_filter_coefs[2][184] = 16'h0000;
	mel_filter_coefs[2][185] = 16'h0000;
	mel_filter_coefs[2][186] = 16'h0000;
	mel_filter_coefs[2][187] = 16'h0000;
	mel_filter_coefs[2][188] = 16'h0000;
	mel_filter_coefs[2][189] = 16'h0000;
	mel_filter_coefs[2][190] = 16'h0000;
	mel_filter_coefs[2][191] = 16'h0000;
	mel_filter_coefs[2][192] = 16'h0000;
	mel_filter_coefs[2][193] = 16'h0000;
	mel_filter_coefs[2][194] = 16'h0000;
	mel_filter_coefs[2][195] = 16'h0000;
	mel_filter_coefs[2][196] = 16'h0000;
	mel_filter_coefs[2][197] = 16'h0000;
	mel_filter_coefs[2][198] = 16'h0000;
	mel_filter_coefs[2][199] = 16'h0000;
	mel_filter_coefs[2][200] = 16'h0000;
	mel_filter_coefs[2][201] = 16'h0000;
	mel_filter_coefs[2][202] = 16'h0000;
	mel_filter_coefs[2][203] = 16'h0000;
	mel_filter_coefs[2][204] = 16'h0000;
	mel_filter_coefs[2][205] = 16'h0000;
	mel_filter_coefs[2][206] = 16'h0000;
	mel_filter_coefs[2][207] = 16'h0000;
	mel_filter_coefs[2][208] = 16'h0000;
	mel_filter_coefs[2][209] = 16'h0000;
	mel_filter_coefs[2][210] = 16'h0000;
	mel_filter_coefs[2][211] = 16'h0000;
	mel_filter_coefs[2][212] = 16'h0000;
	mel_filter_coefs[2][213] = 16'h0000;
	mel_filter_coefs[2][214] = 16'h0000;
	mel_filter_coefs[2][215] = 16'h0000;
	mel_filter_coefs[2][216] = 16'h0000;
	mel_filter_coefs[2][217] = 16'h0000;
	mel_filter_coefs[2][218] = 16'h0000;
	mel_filter_coefs[2][219] = 16'h0000;
	mel_filter_coefs[2][220] = 16'h0000;
	mel_filter_coefs[2][221] = 16'h0000;
	mel_filter_coefs[2][222] = 16'h0000;
	mel_filter_coefs[2][223] = 16'h0000;
	mel_filter_coefs[2][224] = 16'h0000;
	mel_filter_coefs[2][225] = 16'h0000;
	mel_filter_coefs[2][226] = 16'h0000;
	mel_filter_coefs[2][227] = 16'h0000;
	mel_filter_coefs[2][228] = 16'h0000;
	mel_filter_coefs[2][229] = 16'h0000;
	mel_filter_coefs[2][230] = 16'h0000;
	mel_filter_coefs[2][231] = 16'h0000;
	mel_filter_coefs[2][232] = 16'h0000;
	mel_filter_coefs[2][233] = 16'h0000;
	mel_filter_coefs[2][234] = 16'h0000;
	mel_filter_coefs[2][235] = 16'h0000;
	mel_filter_coefs[2][236] = 16'h0000;
	mel_filter_coefs[2][237] = 16'h0000;
	mel_filter_coefs[2][238] = 16'h0000;
	mel_filter_coefs[2][239] = 16'h0000;
	mel_filter_coefs[2][240] = 16'h0000;
	mel_filter_coefs[2][241] = 16'h0000;
	mel_filter_coefs[2][242] = 16'h0000;
	mel_filter_coefs[2][243] = 16'h0000;
	mel_filter_coefs[2][244] = 16'h0000;
	mel_filter_coefs[2][245] = 16'h0000;
	mel_filter_coefs[2][246] = 16'h0000;
	mel_filter_coefs[2][247] = 16'h0000;
	mel_filter_coefs[2][248] = 16'h0000;
	mel_filter_coefs[2][249] = 16'h0000;
	mel_filter_coefs[2][250] = 16'h0000;
	mel_filter_coefs[2][251] = 16'h0000;
	mel_filter_coefs[2][252] = 16'h0000;
	mel_filter_coefs[2][253] = 16'h0000;
	mel_filter_coefs[2][254] = 16'h0000;
	mel_filter_coefs[2][255] = 16'h0000;
	mel_filter_coefs[3][0] = 16'h0000;
	mel_filter_coefs[3][1] = 16'h0000;
	mel_filter_coefs[3][2] = 16'h0000;
	mel_filter_coefs[3][3] = 16'h0000;
	mel_filter_coefs[3][4] = 16'h0000;
	mel_filter_coefs[3][5] = 16'h2447;
	mel_filter_coefs[3][6] = 16'h6F89;
	mel_filter_coefs[3][7] = 16'h48B6;
	mel_filter_coefs[3][8] = 16'h01F1;
	mel_filter_coefs[3][9] = 16'h0000;
	mel_filter_coefs[3][10] = 16'h0000;
	mel_filter_coefs[3][11] = 16'h0000;
	mel_filter_coefs[3][12] = 16'h0000;
	mel_filter_coefs[3][13] = 16'h0000;
	mel_filter_coefs[3][14] = 16'h0000;
	mel_filter_coefs[3][15] = 16'h0000;
	mel_filter_coefs[3][16] = 16'h0000;
	mel_filter_coefs[3][17] = 16'h0000;
	mel_filter_coefs[3][18] = 16'h0000;
	mel_filter_coefs[3][19] = 16'h0000;
	mel_filter_coefs[3][20] = 16'h0000;
	mel_filter_coefs[3][21] = 16'h0000;
	mel_filter_coefs[3][22] = 16'h0000;
	mel_filter_coefs[3][23] = 16'h0000;
	mel_filter_coefs[3][24] = 16'h0000;
	mel_filter_coefs[3][25] = 16'h0000;
	mel_filter_coefs[3][26] = 16'h0000;
	mel_filter_coefs[3][27] = 16'h0000;
	mel_filter_coefs[3][28] = 16'h0000;
	mel_filter_coefs[3][29] = 16'h0000;
	mel_filter_coefs[3][30] = 16'h0000;
	mel_filter_coefs[3][31] = 16'h0000;
	mel_filter_coefs[3][32] = 16'h0000;
	mel_filter_coefs[3][33] = 16'h0000;
	mel_filter_coefs[3][34] = 16'h0000;
	mel_filter_coefs[3][35] = 16'h0000;
	mel_filter_coefs[3][36] = 16'h0000;
	mel_filter_coefs[3][37] = 16'h0000;
	mel_filter_coefs[3][38] = 16'h0000;
	mel_filter_coefs[3][39] = 16'h0000;
	mel_filter_coefs[3][40] = 16'h0000;
	mel_filter_coefs[3][41] = 16'h0000;
	mel_filter_coefs[3][42] = 16'h0000;
	mel_filter_coefs[3][43] = 16'h0000;
	mel_filter_coefs[3][44] = 16'h0000;
	mel_filter_coefs[3][45] = 16'h0000;
	mel_filter_coefs[3][46] = 16'h0000;
	mel_filter_coefs[3][47] = 16'h0000;
	mel_filter_coefs[3][48] = 16'h0000;
	mel_filter_coefs[3][49] = 16'h0000;
	mel_filter_coefs[3][50] = 16'h0000;
	mel_filter_coefs[3][51] = 16'h0000;
	mel_filter_coefs[3][52] = 16'h0000;
	mel_filter_coefs[3][53] = 16'h0000;
	mel_filter_coefs[3][54] = 16'h0000;
	mel_filter_coefs[3][55] = 16'h0000;
	mel_filter_coefs[3][56] = 16'h0000;
	mel_filter_coefs[3][57] = 16'h0000;
	mel_filter_coefs[3][58] = 16'h0000;
	mel_filter_coefs[3][59] = 16'h0000;
	mel_filter_coefs[3][60] = 16'h0000;
	mel_filter_coefs[3][61] = 16'h0000;
	mel_filter_coefs[3][62] = 16'h0000;
	mel_filter_coefs[3][63] = 16'h0000;
	mel_filter_coefs[3][64] = 16'h0000;
	mel_filter_coefs[3][65] = 16'h0000;
	mel_filter_coefs[3][66] = 16'h0000;
	mel_filter_coefs[3][67] = 16'h0000;
	mel_filter_coefs[3][68] = 16'h0000;
	mel_filter_coefs[3][69] = 16'h0000;
	mel_filter_coefs[3][70] = 16'h0000;
	mel_filter_coefs[3][71] = 16'h0000;
	mel_filter_coefs[3][72] = 16'h0000;
	mel_filter_coefs[3][73] = 16'h0000;
	mel_filter_coefs[3][74] = 16'h0000;
	mel_filter_coefs[3][75] = 16'h0000;
	mel_filter_coefs[3][76] = 16'h0000;
	mel_filter_coefs[3][77] = 16'h0000;
	mel_filter_coefs[3][78] = 16'h0000;
	mel_filter_coefs[3][79] = 16'h0000;
	mel_filter_coefs[3][80] = 16'h0000;
	mel_filter_coefs[3][81] = 16'h0000;
	mel_filter_coefs[3][82] = 16'h0000;
	mel_filter_coefs[3][83] = 16'h0000;
	mel_filter_coefs[3][84] = 16'h0000;
	mel_filter_coefs[3][85] = 16'h0000;
	mel_filter_coefs[3][86] = 16'h0000;
	mel_filter_coefs[3][87] = 16'h0000;
	mel_filter_coefs[3][88] = 16'h0000;
	mel_filter_coefs[3][89] = 16'h0000;
	mel_filter_coefs[3][90] = 16'h0000;
	mel_filter_coefs[3][91] = 16'h0000;
	mel_filter_coefs[3][92] = 16'h0000;
	mel_filter_coefs[3][93] = 16'h0000;
	mel_filter_coefs[3][94] = 16'h0000;
	mel_filter_coefs[3][95] = 16'h0000;
	mel_filter_coefs[3][96] = 16'h0000;
	mel_filter_coefs[3][97] = 16'h0000;
	mel_filter_coefs[3][98] = 16'h0000;
	mel_filter_coefs[3][99] = 16'h0000;
	mel_filter_coefs[3][100] = 16'h0000;
	mel_filter_coefs[3][101] = 16'h0000;
	mel_filter_coefs[3][102] = 16'h0000;
	mel_filter_coefs[3][103] = 16'h0000;
	mel_filter_coefs[3][104] = 16'h0000;
	mel_filter_coefs[3][105] = 16'h0000;
	mel_filter_coefs[3][106] = 16'h0000;
	mel_filter_coefs[3][107] = 16'h0000;
	mel_filter_coefs[3][108] = 16'h0000;
	mel_filter_coefs[3][109] = 16'h0000;
	mel_filter_coefs[3][110] = 16'h0000;
	mel_filter_coefs[3][111] = 16'h0000;
	mel_filter_coefs[3][112] = 16'h0000;
	mel_filter_coefs[3][113] = 16'h0000;
	mel_filter_coefs[3][114] = 16'h0000;
	mel_filter_coefs[3][115] = 16'h0000;
	mel_filter_coefs[3][116] = 16'h0000;
	mel_filter_coefs[3][117] = 16'h0000;
	mel_filter_coefs[3][118] = 16'h0000;
	mel_filter_coefs[3][119] = 16'h0000;
	mel_filter_coefs[3][120] = 16'h0000;
	mel_filter_coefs[3][121] = 16'h0000;
	mel_filter_coefs[3][122] = 16'h0000;
	mel_filter_coefs[3][123] = 16'h0000;
	mel_filter_coefs[3][124] = 16'h0000;
	mel_filter_coefs[3][125] = 16'h0000;
	mel_filter_coefs[3][126] = 16'h0000;
	mel_filter_coefs[3][127] = 16'h0000;
	mel_filter_coefs[3][128] = 16'h0000;
	mel_filter_coefs[3][129] = 16'h0000;
	mel_filter_coefs[3][130] = 16'h0000;
	mel_filter_coefs[3][131] = 16'h0000;
	mel_filter_coefs[3][132] = 16'h0000;
	mel_filter_coefs[3][133] = 16'h0000;
	mel_filter_coefs[3][134] = 16'h0000;
	mel_filter_coefs[3][135] = 16'h0000;
	mel_filter_coefs[3][136] = 16'h0000;
	mel_filter_coefs[3][137] = 16'h0000;
	mel_filter_coefs[3][138] = 16'h0000;
	mel_filter_coefs[3][139] = 16'h0000;
	mel_filter_coefs[3][140] = 16'h0000;
	mel_filter_coefs[3][141] = 16'h0000;
	mel_filter_coefs[3][142] = 16'h0000;
	mel_filter_coefs[3][143] = 16'h0000;
	mel_filter_coefs[3][144] = 16'h0000;
	mel_filter_coefs[3][145] = 16'h0000;
	mel_filter_coefs[3][146] = 16'h0000;
	mel_filter_coefs[3][147] = 16'h0000;
	mel_filter_coefs[3][148] = 16'h0000;
	mel_filter_coefs[3][149] = 16'h0000;
	mel_filter_coefs[3][150] = 16'h0000;
	mel_filter_coefs[3][151] = 16'h0000;
	mel_filter_coefs[3][152] = 16'h0000;
	mel_filter_coefs[3][153] = 16'h0000;
	mel_filter_coefs[3][154] = 16'h0000;
	mel_filter_coefs[3][155] = 16'h0000;
	mel_filter_coefs[3][156] = 16'h0000;
	mel_filter_coefs[3][157] = 16'h0000;
	mel_filter_coefs[3][158] = 16'h0000;
	mel_filter_coefs[3][159] = 16'h0000;
	mel_filter_coefs[3][160] = 16'h0000;
	mel_filter_coefs[3][161] = 16'h0000;
	mel_filter_coefs[3][162] = 16'h0000;
	mel_filter_coefs[3][163] = 16'h0000;
	mel_filter_coefs[3][164] = 16'h0000;
	mel_filter_coefs[3][165] = 16'h0000;
	mel_filter_coefs[3][166] = 16'h0000;
	mel_filter_coefs[3][167] = 16'h0000;
	mel_filter_coefs[3][168] = 16'h0000;
	mel_filter_coefs[3][169] = 16'h0000;
	mel_filter_coefs[3][170] = 16'h0000;
	mel_filter_coefs[3][171] = 16'h0000;
	mel_filter_coefs[3][172] = 16'h0000;
	mel_filter_coefs[3][173] = 16'h0000;
	mel_filter_coefs[3][174] = 16'h0000;
	mel_filter_coefs[3][175] = 16'h0000;
	mel_filter_coefs[3][176] = 16'h0000;
	mel_filter_coefs[3][177] = 16'h0000;
	mel_filter_coefs[3][178] = 16'h0000;
	mel_filter_coefs[3][179] = 16'h0000;
	mel_filter_coefs[3][180] = 16'h0000;
	mel_filter_coefs[3][181] = 16'h0000;
	mel_filter_coefs[3][182] = 16'h0000;
	mel_filter_coefs[3][183] = 16'h0000;
	mel_filter_coefs[3][184] = 16'h0000;
	mel_filter_coefs[3][185] = 16'h0000;
	mel_filter_coefs[3][186] = 16'h0000;
	mel_filter_coefs[3][187] = 16'h0000;
	mel_filter_coefs[3][188] = 16'h0000;
	mel_filter_coefs[3][189] = 16'h0000;
	mel_filter_coefs[3][190] = 16'h0000;
	mel_filter_coefs[3][191] = 16'h0000;
	mel_filter_coefs[3][192] = 16'h0000;
	mel_filter_coefs[3][193] = 16'h0000;
	mel_filter_coefs[3][194] = 16'h0000;
	mel_filter_coefs[3][195] = 16'h0000;
	mel_filter_coefs[3][196] = 16'h0000;
	mel_filter_coefs[3][197] = 16'h0000;
	mel_filter_coefs[3][198] = 16'h0000;
	mel_filter_coefs[3][199] = 16'h0000;
	mel_filter_coefs[3][200] = 16'h0000;
	mel_filter_coefs[3][201] = 16'h0000;
	mel_filter_coefs[3][202] = 16'h0000;
	mel_filter_coefs[3][203] = 16'h0000;
	mel_filter_coefs[3][204] = 16'h0000;
	mel_filter_coefs[3][205] = 16'h0000;
	mel_filter_coefs[3][206] = 16'h0000;
	mel_filter_coefs[3][207] = 16'h0000;
	mel_filter_coefs[3][208] = 16'h0000;
	mel_filter_coefs[3][209] = 16'h0000;
	mel_filter_coefs[3][210] = 16'h0000;
	mel_filter_coefs[3][211] = 16'h0000;
	mel_filter_coefs[3][212] = 16'h0000;
	mel_filter_coefs[3][213] = 16'h0000;
	mel_filter_coefs[3][214] = 16'h0000;
	mel_filter_coefs[3][215] = 16'h0000;
	mel_filter_coefs[3][216] = 16'h0000;
	mel_filter_coefs[3][217] = 16'h0000;
	mel_filter_coefs[3][218] = 16'h0000;
	mel_filter_coefs[3][219] = 16'h0000;
	mel_filter_coefs[3][220] = 16'h0000;
	mel_filter_coefs[3][221] = 16'h0000;
	mel_filter_coefs[3][222] = 16'h0000;
	mel_filter_coefs[3][223] = 16'h0000;
	mel_filter_coefs[3][224] = 16'h0000;
	mel_filter_coefs[3][225] = 16'h0000;
	mel_filter_coefs[3][226] = 16'h0000;
	mel_filter_coefs[3][227] = 16'h0000;
	mel_filter_coefs[3][228] = 16'h0000;
	mel_filter_coefs[3][229] = 16'h0000;
	mel_filter_coefs[3][230] = 16'h0000;
	mel_filter_coefs[3][231] = 16'h0000;
	mel_filter_coefs[3][232] = 16'h0000;
	mel_filter_coefs[3][233] = 16'h0000;
	mel_filter_coefs[3][234] = 16'h0000;
	mel_filter_coefs[3][235] = 16'h0000;
	mel_filter_coefs[3][236] = 16'h0000;
	mel_filter_coefs[3][237] = 16'h0000;
	mel_filter_coefs[3][238] = 16'h0000;
	mel_filter_coefs[3][239] = 16'h0000;
	mel_filter_coefs[3][240] = 16'h0000;
	mel_filter_coefs[3][241] = 16'h0000;
	mel_filter_coefs[3][242] = 16'h0000;
	mel_filter_coefs[3][243] = 16'h0000;
	mel_filter_coefs[3][244] = 16'h0000;
	mel_filter_coefs[3][245] = 16'h0000;
	mel_filter_coefs[3][246] = 16'h0000;
	mel_filter_coefs[3][247] = 16'h0000;
	mel_filter_coefs[3][248] = 16'h0000;
	mel_filter_coefs[3][249] = 16'h0000;
	mel_filter_coefs[3][250] = 16'h0000;
	mel_filter_coefs[3][251] = 16'h0000;
	mel_filter_coefs[3][252] = 16'h0000;
	mel_filter_coefs[3][253] = 16'h0000;
	mel_filter_coefs[3][254] = 16'h0000;
	mel_filter_coefs[3][255] = 16'h0000;
	mel_filter_coefs[4][0] = 16'h0000;
	mel_filter_coefs[4][1] = 16'h0000;
	mel_filter_coefs[4][2] = 16'h0000;
	mel_filter_coefs[4][3] = 16'h0000;
	mel_filter_coefs[4][4] = 16'h0000;
	mel_filter_coefs[4][5] = 16'h0000;
	mel_filter_coefs[4][6] = 16'h0000;
	mel_filter_coefs[4][7] = 16'h374A;
	mel_filter_coefs[4][8] = 16'h7E0F;
	mel_filter_coefs[4][9] = 16'h3F45;
	mel_filter_coefs[4][10] = 16'h0000;
	mel_filter_coefs[4][11] = 16'h0000;
	mel_filter_coefs[4][12] = 16'h0000;
	mel_filter_coefs[4][13] = 16'h0000;
	mel_filter_coefs[4][14] = 16'h0000;
	mel_filter_coefs[4][15] = 16'h0000;
	mel_filter_coefs[4][16] = 16'h0000;
	mel_filter_coefs[4][17] = 16'h0000;
	mel_filter_coefs[4][18] = 16'h0000;
	mel_filter_coefs[4][19] = 16'h0000;
	mel_filter_coefs[4][20] = 16'h0000;
	mel_filter_coefs[4][21] = 16'h0000;
	mel_filter_coefs[4][22] = 16'h0000;
	mel_filter_coefs[4][23] = 16'h0000;
	mel_filter_coefs[4][24] = 16'h0000;
	mel_filter_coefs[4][25] = 16'h0000;
	mel_filter_coefs[4][26] = 16'h0000;
	mel_filter_coefs[4][27] = 16'h0000;
	mel_filter_coefs[4][28] = 16'h0000;
	mel_filter_coefs[4][29] = 16'h0000;
	mel_filter_coefs[4][30] = 16'h0000;
	mel_filter_coefs[4][31] = 16'h0000;
	mel_filter_coefs[4][32] = 16'h0000;
	mel_filter_coefs[4][33] = 16'h0000;
	mel_filter_coefs[4][34] = 16'h0000;
	mel_filter_coefs[4][35] = 16'h0000;
	mel_filter_coefs[4][36] = 16'h0000;
	mel_filter_coefs[4][37] = 16'h0000;
	mel_filter_coefs[4][38] = 16'h0000;
	mel_filter_coefs[4][39] = 16'h0000;
	mel_filter_coefs[4][40] = 16'h0000;
	mel_filter_coefs[4][41] = 16'h0000;
	mel_filter_coefs[4][42] = 16'h0000;
	mel_filter_coefs[4][43] = 16'h0000;
	mel_filter_coefs[4][44] = 16'h0000;
	mel_filter_coefs[4][45] = 16'h0000;
	mel_filter_coefs[4][46] = 16'h0000;
	mel_filter_coefs[4][47] = 16'h0000;
	mel_filter_coefs[4][48] = 16'h0000;
	mel_filter_coefs[4][49] = 16'h0000;
	mel_filter_coefs[4][50] = 16'h0000;
	mel_filter_coefs[4][51] = 16'h0000;
	mel_filter_coefs[4][52] = 16'h0000;
	mel_filter_coefs[4][53] = 16'h0000;
	mel_filter_coefs[4][54] = 16'h0000;
	mel_filter_coefs[4][55] = 16'h0000;
	mel_filter_coefs[4][56] = 16'h0000;
	mel_filter_coefs[4][57] = 16'h0000;
	mel_filter_coefs[4][58] = 16'h0000;
	mel_filter_coefs[4][59] = 16'h0000;
	mel_filter_coefs[4][60] = 16'h0000;
	mel_filter_coefs[4][61] = 16'h0000;
	mel_filter_coefs[4][62] = 16'h0000;
	mel_filter_coefs[4][63] = 16'h0000;
	mel_filter_coefs[4][64] = 16'h0000;
	mel_filter_coefs[4][65] = 16'h0000;
	mel_filter_coefs[4][66] = 16'h0000;
	mel_filter_coefs[4][67] = 16'h0000;
	mel_filter_coefs[4][68] = 16'h0000;
	mel_filter_coefs[4][69] = 16'h0000;
	mel_filter_coefs[4][70] = 16'h0000;
	mel_filter_coefs[4][71] = 16'h0000;
	mel_filter_coefs[4][72] = 16'h0000;
	mel_filter_coefs[4][73] = 16'h0000;
	mel_filter_coefs[4][74] = 16'h0000;
	mel_filter_coefs[4][75] = 16'h0000;
	mel_filter_coefs[4][76] = 16'h0000;
	mel_filter_coefs[4][77] = 16'h0000;
	mel_filter_coefs[4][78] = 16'h0000;
	mel_filter_coefs[4][79] = 16'h0000;
	mel_filter_coefs[4][80] = 16'h0000;
	mel_filter_coefs[4][81] = 16'h0000;
	mel_filter_coefs[4][82] = 16'h0000;
	mel_filter_coefs[4][83] = 16'h0000;
	mel_filter_coefs[4][84] = 16'h0000;
	mel_filter_coefs[4][85] = 16'h0000;
	mel_filter_coefs[4][86] = 16'h0000;
	mel_filter_coefs[4][87] = 16'h0000;
	mel_filter_coefs[4][88] = 16'h0000;
	mel_filter_coefs[4][89] = 16'h0000;
	mel_filter_coefs[4][90] = 16'h0000;
	mel_filter_coefs[4][91] = 16'h0000;
	mel_filter_coefs[4][92] = 16'h0000;
	mel_filter_coefs[4][93] = 16'h0000;
	mel_filter_coefs[4][94] = 16'h0000;
	mel_filter_coefs[4][95] = 16'h0000;
	mel_filter_coefs[4][96] = 16'h0000;
	mel_filter_coefs[4][97] = 16'h0000;
	mel_filter_coefs[4][98] = 16'h0000;
	mel_filter_coefs[4][99] = 16'h0000;
	mel_filter_coefs[4][100] = 16'h0000;
	mel_filter_coefs[4][101] = 16'h0000;
	mel_filter_coefs[4][102] = 16'h0000;
	mel_filter_coefs[4][103] = 16'h0000;
	mel_filter_coefs[4][104] = 16'h0000;
	mel_filter_coefs[4][105] = 16'h0000;
	mel_filter_coefs[4][106] = 16'h0000;
	mel_filter_coefs[4][107] = 16'h0000;
	mel_filter_coefs[4][108] = 16'h0000;
	mel_filter_coefs[4][109] = 16'h0000;
	mel_filter_coefs[4][110] = 16'h0000;
	mel_filter_coefs[4][111] = 16'h0000;
	mel_filter_coefs[4][112] = 16'h0000;
	mel_filter_coefs[4][113] = 16'h0000;
	mel_filter_coefs[4][114] = 16'h0000;
	mel_filter_coefs[4][115] = 16'h0000;
	mel_filter_coefs[4][116] = 16'h0000;
	mel_filter_coefs[4][117] = 16'h0000;
	mel_filter_coefs[4][118] = 16'h0000;
	mel_filter_coefs[4][119] = 16'h0000;
	mel_filter_coefs[4][120] = 16'h0000;
	mel_filter_coefs[4][121] = 16'h0000;
	mel_filter_coefs[4][122] = 16'h0000;
	mel_filter_coefs[4][123] = 16'h0000;
	mel_filter_coefs[4][124] = 16'h0000;
	mel_filter_coefs[4][125] = 16'h0000;
	mel_filter_coefs[4][126] = 16'h0000;
	mel_filter_coefs[4][127] = 16'h0000;
	mel_filter_coefs[4][128] = 16'h0000;
	mel_filter_coefs[4][129] = 16'h0000;
	mel_filter_coefs[4][130] = 16'h0000;
	mel_filter_coefs[4][131] = 16'h0000;
	mel_filter_coefs[4][132] = 16'h0000;
	mel_filter_coefs[4][133] = 16'h0000;
	mel_filter_coefs[4][134] = 16'h0000;
	mel_filter_coefs[4][135] = 16'h0000;
	mel_filter_coefs[4][136] = 16'h0000;
	mel_filter_coefs[4][137] = 16'h0000;
	mel_filter_coefs[4][138] = 16'h0000;
	mel_filter_coefs[4][139] = 16'h0000;
	mel_filter_coefs[4][140] = 16'h0000;
	mel_filter_coefs[4][141] = 16'h0000;
	mel_filter_coefs[4][142] = 16'h0000;
	mel_filter_coefs[4][143] = 16'h0000;
	mel_filter_coefs[4][144] = 16'h0000;
	mel_filter_coefs[4][145] = 16'h0000;
	mel_filter_coefs[4][146] = 16'h0000;
	mel_filter_coefs[4][147] = 16'h0000;
	mel_filter_coefs[4][148] = 16'h0000;
	mel_filter_coefs[4][149] = 16'h0000;
	mel_filter_coefs[4][150] = 16'h0000;
	mel_filter_coefs[4][151] = 16'h0000;
	mel_filter_coefs[4][152] = 16'h0000;
	mel_filter_coefs[4][153] = 16'h0000;
	mel_filter_coefs[4][154] = 16'h0000;
	mel_filter_coefs[4][155] = 16'h0000;
	mel_filter_coefs[4][156] = 16'h0000;
	mel_filter_coefs[4][157] = 16'h0000;
	mel_filter_coefs[4][158] = 16'h0000;
	mel_filter_coefs[4][159] = 16'h0000;
	mel_filter_coefs[4][160] = 16'h0000;
	mel_filter_coefs[4][161] = 16'h0000;
	mel_filter_coefs[4][162] = 16'h0000;
	mel_filter_coefs[4][163] = 16'h0000;
	mel_filter_coefs[4][164] = 16'h0000;
	mel_filter_coefs[4][165] = 16'h0000;
	mel_filter_coefs[4][166] = 16'h0000;
	mel_filter_coefs[4][167] = 16'h0000;
	mel_filter_coefs[4][168] = 16'h0000;
	mel_filter_coefs[4][169] = 16'h0000;
	mel_filter_coefs[4][170] = 16'h0000;
	mel_filter_coefs[4][171] = 16'h0000;
	mel_filter_coefs[4][172] = 16'h0000;
	mel_filter_coefs[4][173] = 16'h0000;
	mel_filter_coefs[4][174] = 16'h0000;
	mel_filter_coefs[4][175] = 16'h0000;
	mel_filter_coefs[4][176] = 16'h0000;
	mel_filter_coefs[4][177] = 16'h0000;
	mel_filter_coefs[4][178] = 16'h0000;
	mel_filter_coefs[4][179] = 16'h0000;
	mel_filter_coefs[4][180] = 16'h0000;
	mel_filter_coefs[4][181] = 16'h0000;
	mel_filter_coefs[4][182] = 16'h0000;
	mel_filter_coefs[4][183] = 16'h0000;
	mel_filter_coefs[4][184] = 16'h0000;
	mel_filter_coefs[4][185] = 16'h0000;
	mel_filter_coefs[4][186] = 16'h0000;
	mel_filter_coefs[4][187] = 16'h0000;
	mel_filter_coefs[4][188] = 16'h0000;
	mel_filter_coefs[4][189] = 16'h0000;
	mel_filter_coefs[4][190] = 16'h0000;
	mel_filter_coefs[4][191] = 16'h0000;
	mel_filter_coefs[4][192] = 16'h0000;
	mel_filter_coefs[4][193] = 16'h0000;
	mel_filter_coefs[4][194] = 16'h0000;
	mel_filter_coefs[4][195] = 16'h0000;
	mel_filter_coefs[4][196] = 16'h0000;
	mel_filter_coefs[4][197] = 16'h0000;
	mel_filter_coefs[4][198] = 16'h0000;
	mel_filter_coefs[4][199] = 16'h0000;
	mel_filter_coefs[4][200] = 16'h0000;
	mel_filter_coefs[4][201] = 16'h0000;
	mel_filter_coefs[4][202] = 16'h0000;
	mel_filter_coefs[4][203] = 16'h0000;
	mel_filter_coefs[4][204] = 16'h0000;
	mel_filter_coefs[4][205] = 16'h0000;
	mel_filter_coefs[4][206] = 16'h0000;
	mel_filter_coefs[4][207] = 16'h0000;
	mel_filter_coefs[4][208] = 16'h0000;
	mel_filter_coefs[4][209] = 16'h0000;
	mel_filter_coefs[4][210] = 16'h0000;
	mel_filter_coefs[4][211] = 16'h0000;
	mel_filter_coefs[4][212] = 16'h0000;
	mel_filter_coefs[4][213] = 16'h0000;
	mel_filter_coefs[4][214] = 16'h0000;
	mel_filter_coefs[4][215] = 16'h0000;
	mel_filter_coefs[4][216] = 16'h0000;
	mel_filter_coefs[4][217] = 16'h0000;
	mel_filter_coefs[4][218] = 16'h0000;
	mel_filter_coefs[4][219] = 16'h0000;
	mel_filter_coefs[4][220] = 16'h0000;
	mel_filter_coefs[4][221] = 16'h0000;
	mel_filter_coefs[4][222] = 16'h0000;
	mel_filter_coefs[4][223] = 16'h0000;
	mel_filter_coefs[4][224] = 16'h0000;
	mel_filter_coefs[4][225] = 16'h0000;
	mel_filter_coefs[4][226] = 16'h0000;
	mel_filter_coefs[4][227] = 16'h0000;
	mel_filter_coefs[4][228] = 16'h0000;
	mel_filter_coefs[4][229] = 16'h0000;
	mel_filter_coefs[4][230] = 16'h0000;
	mel_filter_coefs[4][231] = 16'h0000;
	mel_filter_coefs[4][232] = 16'h0000;
	mel_filter_coefs[4][233] = 16'h0000;
	mel_filter_coefs[4][234] = 16'h0000;
	mel_filter_coefs[4][235] = 16'h0000;
	mel_filter_coefs[4][236] = 16'h0000;
	mel_filter_coefs[4][237] = 16'h0000;
	mel_filter_coefs[4][238] = 16'h0000;
	mel_filter_coefs[4][239] = 16'h0000;
	mel_filter_coefs[4][240] = 16'h0000;
	mel_filter_coefs[4][241] = 16'h0000;
	mel_filter_coefs[4][242] = 16'h0000;
	mel_filter_coefs[4][243] = 16'h0000;
	mel_filter_coefs[4][244] = 16'h0000;
	mel_filter_coefs[4][245] = 16'h0000;
	mel_filter_coefs[4][246] = 16'h0000;
	mel_filter_coefs[4][247] = 16'h0000;
	mel_filter_coefs[4][248] = 16'h0000;
	mel_filter_coefs[4][249] = 16'h0000;
	mel_filter_coefs[4][250] = 16'h0000;
	mel_filter_coefs[4][251] = 16'h0000;
	mel_filter_coefs[4][252] = 16'h0000;
	mel_filter_coefs[4][253] = 16'h0000;
	mel_filter_coefs[4][254] = 16'h0000;
	mel_filter_coefs[4][255] = 16'h0000;
	mel_filter_coefs[5][0] = 16'h0000;
	mel_filter_coefs[5][1] = 16'h0000;
	mel_filter_coefs[5][2] = 16'h0000;
	mel_filter_coefs[5][3] = 16'h0000;
	mel_filter_coefs[5][4] = 16'h0000;
	mel_filter_coefs[5][5] = 16'h0000;
	mel_filter_coefs[5][6] = 16'h0000;
	mel_filter_coefs[5][7] = 16'h0000;
	mel_filter_coefs[5][8] = 16'h0000;
	mel_filter_coefs[5][9] = 16'h40BB;
	mel_filter_coefs[5][10] = 16'h7CEA;
	mel_filter_coefs[5][11] = 16'h3E54;
	mel_filter_coefs[5][12] = 16'h0000;
	mel_filter_coefs[5][13] = 16'h0000;
	mel_filter_coefs[5][14] = 16'h0000;
	mel_filter_coefs[5][15] = 16'h0000;
	mel_filter_coefs[5][16] = 16'h0000;
	mel_filter_coefs[5][17] = 16'h0000;
	mel_filter_coefs[5][18] = 16'h0000;
	mel_filter_coefs[5][19] = 16'h0000;
	mel_filter_coefs[5][20] = 16'h0000;
	mel_filter_coefs[5][21] = 16'h0000;
	mel_filter_coefs[5][22] = 16'h0000;
	mel_filter_coefs[5][23] = 16'h0000;
	mel_filter_coefs[5][24] = 16'h0000;
	mel_filter_coefs[5][25] = 16'h0000;
	mel_filter_coefs[5][26] = 16'h0000;
	mel_filter_coefs[5][27] = 16'h0000;
	mel_filter_coefs[5][28] = 16'h0000;
	mel_filter_coefs[5][29] = 16'h0000;
	mel_filter_coefs[5][30] = 16'h0000;
	mel_filter_coefs[5][31] = 16'h0000;
	mel_filter_coefs[5][32] = 16'h0000;
	mel_filter_coefs[5][33] = 16'h0000;
	mel_filter_coefs[5][34] = 16'h0000;
	mel_filter_coefs[5][35] = 16'h0000;
	mel_filter_coefs[5][36] = 16'h0000;
	mel_filter_coefs[5][37] = 16'h0000;
	mel_filter_coefs[5][38] = 16'h0000;
	mel_filter_coefs[5][39] = 16'h0000;
	mel_filter_coefs[5][40] = 16'h0000;
	mel_filter_coefs[5][41] = 16'h0000;
	mel_filter_coefs[5][42] = 16'h0000;
	mel_filter_coefs[5][43] = 16'h0000;
	mel_filter_coefs[5][44] = 16'h0000;
	mel_filter_coefs[5][45] = 16'h0000;
	mel_filter_coefs[5][46] = 16'h0000;
	mel_filter_coefs[5][47] = 16'h0000;
	mel_filter_coefs[5][48] = 16'h0000;
	mel_filter_coefs[5][49] = 16'h0000;
	mel_filter_coefs[5][50] = 16'h0000;
	mel_filter_coefs[5][51] = 16'h0000;
	mel_filter_coefs[5][52] = 16'h0000;
	mel_filter_coefs[5][53] = 16'h0000;
	mel_filter_coefs[5][54] = 16'h0000;
	mel_filter_coefs[5][55] = 16'h0000;
	mel_filter_coefs[5][56] = 16'h0000;
	mel_filter_coefs[5][57] = 16'h0000;
	mel_filter_coefs[5][58] = 16'h0000;
	mel_filter_coefs[5][59] = 16'h0000;
	mel_filter_coefs[5][60] = 16'h0000;
	mel_filter_coefs[5][61] = 16'h0000;
	mel_filter_coefs[5][62] = 16'h0000;
	mel_filter_coefs[5][63] = 16'h0000;
	mel_filter_coefs[5][64] = 16'h0000;
	mel_filter_coefs[5][65] = 16'h0000;
	mel_filter_coefs[5][66] = 16'h0000;
	mel_filter_coefs[5][67] = 16'h0000;
	mel_filter_coefs[5][68] = 16'h0000;
	mel_filter_coefs[5][69] = 16'h0000;
	mel_filter_coefs[5][70] = 16'h0000;
	mel_filter_coefs[5][71] = 16'h0000;
	mel_filter_coefs[5][72] = 16'h0000;
	mel_filter_coefs[5][73] = 16'h0000;
	mel_filter_coefs[5][74] = 16'h0000;
	mel_filter_coefs[5][75] = 16'h0000;
	mel_filter_coefs[5][76] = 16'h0000;
	mel_filter_coefs[5][77] = 16'h0000;
	mel_filter_coefs[5][78] = 16'h0000;
	mel_filter_coefs[5][79] = 16'h0000;
	mel_filter_coefs[5][80] = 16'h0000;
	mel_filter_coefs[5][81] = 16'h0000;
	mel_filter_coefs[5][82] = 16'h0000;
	mel_filter_coefs[5][83] = 16'h0000;
	mel_filter_coefs[5][84] = 16'h0000;
	mel_filter_coefs[5][85] = 16'h0000;
	mel_filter_coefs[5][86] = 16'h0000;
	mel_filter_coefs[5][87] = 16'h0000;
	mel_filter_coefs[5][88] = 16'h0000;
	mel_filter_coefs[5][89] = 16'h0000;
	mel_filter_coefs[5][90] = 16'h0000;
	mel_filter_coefs[5][91] = 16'h0000;
	mel_filter_coefs[5][92] = 16'h0000;
	mel_filter_coefs[5][93] = 16'h0000;
	mel_filter_coefs[5][94] = 16'h0000;
	mel_filter_coefs[5][95] = 16'h0000;
	mel_filter_coefs[5][96] = 16'h0000;
	mel_filter_coefs[5][97] = 16'h0000;
	mel_filter_coefs[5][98] = 16'h0000;
	mel_filter_coefs[5][99] = 16'h0000;
	mel_filter_coefs[5][100] = 16'h0000;
	mel_filter_coefs[5][101] = 16'h0000;
	mel_filter_coefs[5][102] = 16'h0000;
	mel_filter_coefs[5][103] = 16'h0000;
	mel_filter_coefs[5][104] = 16'h0000;
	mel_filter_coefs[5][105] = 16'h0000;
	mel_filter_coefs[5][106] = 16'h0000;
	mel_filter_coefs[5][107] = 16'h0000;
	mel_filter_coefs[5][108] = 16'h0000;
	mel_filter_coefs[5][109] = 16'h0000;
	mel_filter_coefs[5][110] = 16'h0000;
	mel_filter_coefs[5][111] = 16'h0000;
	mel_filter_coefs[5][112] = 16'h0000;
	mel_filter_coefs[5][113] = 16'h0000;
	mel_filter_coefs[5][114] = 16'h0000;
	mel_filter_coefs[5][115] = 16'h0000;
	mel_filter_coefs[5][116] = 16'h0000;
	mel_filter_coefs[5][117] = 16'h0000;
	mel_filter_coefs[5][118] = 16'h0000;
	mel_filter_coefs[5][119] = 16'h0000;
	mel_filter_coefs[5][120] = 16'h0000;
	mel_filter_coefs[5][121] = 16'h0000;
	mel_filter_coefs[5][122] = 16'h0000;
	mel_filter_coefs[5][123] = 16'h0000;
	mel_filter_coefs[5][124] = 16'h0000;
	mel_filter_coefs[5][125] = 16'h0000;
	mel_filter_coefs[5][126] = 16'h0000;
	mel_filter_coefs[5][127] = 16'h0000;
	mel_filter_coefs[5][128] = 16'h0000;
	mel_filter_coefs[5][129] = 16'h0000;
	mel_filter_coefs[5][130] = 16'h0000;
	mel_filter_coefs[5][131] = 16'h0000;
	mel_filter_coefs[5][132] = 16'h0000;
	mel_filter_coefs[5][133] = 16'h0000;
	mel_filter_coefs[5][134] = 16'h0000;
	mel_filter_coefs[5][135] = 16'h0000;
	mel_filter_coefs[5][136] = 16'h0000;
	mel_filter_coefs[5][137] = 16'h0000;
	mel_filter_coefs[5][138] = 16'h0000;
	mel_filter_coefs[5][139] = 16'h0000;
	mel_filter_coefs[5][140] = 16'h0000;
	mel_filter_coefs[5][141] = 16'h0000;
	mel_filter_coefs[5][142] = 16'h0000;
	mel_filter_coefs[5][143] = 16'h0000;
	mel_filter_coefs[5][144] = 16'h0000;
	mel_filter_coefs[5][145] = 16'h0000;
	mel_filter_coefs[5][146] = 16'h0000;
	mel_filter_coefs[5][147] = 16'h0000;
	mel_filter_coefs[5][148] = 16'h0000;
	mel_filter_coefs[5][149] = 16'h0000;
	mel_filter_coefs[5][150] = 16'h0000;
	mel_filter_coefs[5][151] = 16'h0000;
	mel_filter_coefs[5][152] = 16'h0000;
	mel_filter_coefs[5][153] = 16'h0000;
	mel_filter_coefs[5][154] = 16'h0000;
	mel_filter_coefs[5][155] = 16'h0000;
	mel_filter_coefs[5][156] = 16'h0000;
	mel_filter_coefs[5][157] = 16'h0000;
	mel_filter_coefs[5][158] = 16'h0000;
	mel_filter_coefs[5][159] = 16'h0000;
	mel_filter_coefs[5][160] = 16'h0000;
	mel_filter_coefs[5][161] = 16'h0000;
	mel_filter_coefs[5][162] = 16'h0000;
	mel_filter_coefs[5][163] = 16'h0000;
	mel_filter_coefs[5][164] = 16'h0000;
	mel_filter_coefs[5][165] = 16'h0000;
	mel_filter_coefs[5][166] = 16'h0000;
	mel_filter_coefs[5][167] = 16'h0000;
	mel_filter_coefs[5][168] = 16'h0000;
	mel_filter_coefs[5][169] = 16'h0000;
	mel_filter_coefs[5][170] = 16'h0000;
	mel_filter_coefs[5][171] = 16'h0000;
	mel_filter_coefs[5][172] = 16'h0000;
	mel_filter_coefs[5][173] = 16'h0000;
	mel_filter_coefs[5][174] = 16'h0000;
	mel_filter_coefs[5][175] = 16'h0000;
	mel_filter_coefs[5][176] = 16'h0000;
	mel_filter_coefs[5][177] = 16'h0000;
	mel_filter_coefs[5][178] = 16'h0000;
	mel_filter_coefs[5][179] = 16'h0000;
	mel_filter_coefs[5][180] = 16'h0000;
	mel_filter_coefs[5][181] = 16'h0000;
	mel_filter_coefs[5][182] = 16'h0000;
	mel_filter_coefs[5][183] = 16'h0000;
	mel_filter_coefs[5][184] = 16'h0000;
	mel_filter_coefs[5][185] = 16'h0000;
	mel_filter_coefs[5][186] = 16'h0000;
	mel_filter_coefs[5][187] = 16'h0000;
	mel_filter_coefs[5][188] = 16'h0000;
	mel_filter_coefs[5][189] = 16'h0000;
	mel_filter_coefs[5][190] = 16'h0000;
	mel_filter_coefs[5][191] = 16'h0000;
	mel_filter_coefs[5][192] = 16'h0000;
	mel_filter_coefs[5][193] = 16'h0000;
	mel_filter_coefs[5][194] = 16'h0000;
	mel_filter_coefs[5][195] = 16'h0000;
	mel_filter_coefs[5][196] = 16'h0000;
	mel_filter_coefs[5][197] = 16'h0000;
	mel_filter_coefs[5][198] = 16'h0000;
	mel_filter_coefs[5][199] = 16'h0000;
	mel_filter_coefs[5][200] = 16'h0000;
	mel_filter_coefs[5][201] = 16'h0000;
	mel_filter_coefs[5][202] = 16'h0000;
	mel_filter_coefs[5][203] = 16'h0000;
	mel_filter_coefs[5][204] = 16'h0000;
	mel_filter_coefs[5][205] = 16'h0000;
	mel_filter_coefs[5][206] = 16'h0000;
	mel_filter_coefs[5][207] = 16'h0000;
	mel_filter_coefs[5][208] = 16'h0000;
	mel_filter_coefs[5][209] = 16'h0000;
	mel_filter_coefs[5][210] = 16'h0000;
	mel_filter_coefs[5][211] = 16'h0000;
	mel_filter_coefs[5][212] = 16'h0000;
	mel_filter_coefs[5][213] = 16'h0000;
	mel_filter_coefs[5][214] = 16'h0000;
	mel_filter_coefs[5][215] = 16'h0000;
	mel_filter_coefs[5][216] = 16'h0000;
	mel_filter_coefs[5][217] = 16'h0000;
	mel_filter_coefs[5][218] = 16'h0000;
	mel_filter_coefs[5][219] = 16'h0000;
	mel_filter_coefs[5][220] = 16'h0000;
	mel_filter_coefs[5][221] = 16'h0000;
	mel_filter_coefs[5][222] = 16'h0000;
	mel_filter_coefs[5][223] = 16'h0000;
	mel_filter_coefs[5][224] = 16'h0000;
	mel_filter_coefs[5][225] = 16'h0000;
	mel_filter_coefs[5][226] = 16'h0000;
	mel_filter_coefs[5][227] = 16'h0000;
	mel_filter_coefs[5][228] = 16'h0000;
	mel_filter_coefs[5][229] = 16'h0000;
	mel_filter_coefs[5][230] = 16'h0000;
	mel_filter_coefs[5][231] = 16'h0000;
	mel_filter_coefs[5][232] = 16'h0000;
	mel_filter_coefs[5][233] = 16'h0000;
	mel_filter_coefs[5][234] = 16'h0000;
	mel_filter_coefs[5][235] = 16'h0000;
	mel_filter_coefs[5][236] = 16'h0000;
	mel_filter_coefs[5][237] = 16'h0000;
	mel_filter_coefs[5][238] = 16'h0000;
	mel_filter_coefs[5][239] = 16'h0000;
	mel_filter_coefs[5][240] = 16'h0000;
	mel_filter_coefs[5][241] = 16'h0000;
	mel_filter_coefs[5][242] = 16'h0000;
	mel_filter_coefs[5][243] = 16'h0000;
	mel_filter_coefs[5][244] = 16'h0000;
	mel_filter_coefs[5][245] = 16'h0000;
	mel_filter_coefs[5][246] = 16'h0000;
	mel_filter_coefs[5][247] = 16'h0000;
	mel_filter_coefs[5][248] = 16'h0000;
	mel_filter_coefs[5][249] = 16'h0000;
	mel_filter_coefs[5][250] = 16'h0000;
	mel_filter_coefs[5][251] = 16'h0000;
	mel_filter_coefs[5][252] = 16'h0000;
	mel_filter_coefs[5][253] = 16'h0000;
	mel_filter_coefs[5][254] = 16'h0000;
	mel_filter_coefs[5][255] = 16'h0000;
	mel_filter_coefs[6][0] = 16'h0000;
	mel_filter_coefs[6][1] = 16'h0000;
	mel_filter_coefs[6][2] = 16'h0000;
	mel_filter_coefs[6][3] = 16'h0000;
	mel_filter_coefs[6][4] = 16'h0000;
	mel_filter_coefs[6][5] = 16'h0000;
	mel_filter_coefs[6][6] = 16'h0000;
	mel_filter_coefs[6][7] = 16'h0000;
	mel_filter_coefs[6][8] = 16'h0000;
	mel_filter_coefs[6][9] = 16'h0000;
	mel_filter_coefs[6][10] = 16'h0316;
	mel_filter_coefs[6][11] = 16'h41AC;
	mel_filter_coefs[6][12] = 16'h7FC2;
	mel_filter_coefs[6][13] = 16'h44E8;
	mel_filter_coefs[6][14] = 16'h0A0D;
	mel_filter_coefs[6][15] = 16'h0000;
	mel_filter_coefs[6][16] = 16'h0000;
	mel_filter_coefs[6][17] = 16'h0000;
	mel_filter_coefs[6][18] = 16'h0000;
	mel_filter_coefs[6][19] = 16'h0000;
	mel_filter_coefs[6][20] = 16'h0000;
	mel_filter_coefs[6][21] = 16'h0000;
	mel_filter_coefs[6][22] = 16'h0000;
	mel_filter_coefs[6][23] = 16'h0000;
	mel_filter_coefs[6][24] = 16'h0000;
	mel_filter_coefs[6][25] = 16'h0000;
	mel_filter_coefs[6][26] = 16'h0000;
	mel_filter_coefs[6][27] = 16'h0000;
	mel_filter_coefs[6][28] = 16'h0000;
	mel_filter_coefs[6][29] = 16'h0000;
	mel_filter_coefs[6][30] = 16'h0000;
	mel_filter_coefs[6][31] = 16'h0000;
	mel_filter_coefs[6][32] = 16'h0000;
	mel_filter_coefs[6][33] = 16'h0000;
	mel_filter_coefs[6][34] = 16'h0000;
	mel_filter_coefs[6][35] = 16'h0000;
	mel_filter_coefs[6][36] = 16'h0000;
	mel_filter_coefs[6][37] = 16'h0000;
	mel_filter_coefs[6][38] = 16'h0000;
	mel_filter_coefs[6][39] = 16'h0000;
	mel_filter_coefs[6][40] = 16'h0000;
	mel_filter_coefs[6][41] = 16'h0000;
	mel_filter_coefs[6][42] = 16'h0000;
	mel_filter_coefs[6][43] = 16'h0000;
	mel_filter_coefs[6][44] = 16'h0000;
	mel_filter_coefs[6][45] = 16'h0000;
	mel_filter_coefs[6][46] = 16'h0000;
	mel_filter_coefs[6][47] = 16'h0000;
	mel_filter_coefs[6][48] = 16'h0000;
	mel_filter_coefs[6][49] = 16'h0000;
	mel_filter_coefs[6][50] = 16'h0000;
	mel_filter_coefs[6][51] = 16'h0000;
	mel_filter_coefs[6][52] = 16'h0000;
	mel_filter_coefs[6][53] = 16'h0000;
	mel_filter_coefs[6][54] = 16'h0000;
	mel_filter_coefs[6][55] = 16'h0000;
	mel_filter_coefs[6][56] = 16'h0000;
	mel_filter_coefs[6][57] = 16'h0000;
	mel_filter_coefs[6][58] = 16'h0000;
	mel_filter_coefs[6][59] = 16'h0000;
	mel_filter_coefs[6][60] = 16'h0000;
	mel_filter_coefs[6][61] = 16'h0000;
	mel_filter_coefs[6][62] = 16'h0000;
	mel_filter_coefs[6][63] = 16'h0000;
	mel_filter_coefs[6][64] = 16'h0000;
	mel_filter_coefs[6][65] = 16'h0000;
	mel_filter_coefs[6][66] = 16'h0000;
	mel_filter_coefs[6][67] = 16'h0000;
	mel_filter_coefs[6][68] = 16'h0000;
	mel_filter_coefs[6][69] = 16'h0000;
	mel_filter_coefs[6][70] = 16'h0000;
	mel_filter_coefs[6][71] = 16'h0000;
	mel_filter_coefs[6][72] = 16'h0000;
	mel_filter_coefs[6][73] = 16'h0000;
	mel_filter_coefs[6][74] = 16'h0000;
	mel_filter_coefs[6][75] = 16'h0000;
	mel_filter_coefs[6][76] = 16'h0000;
	mel_filter_coefs[6][77] = 16'h0000;
	mel_filter_coefs[6][78] = 16'h0000;
	mel_filter_coefs[6][79] = 16'h0000;
	mel_filter_coefs[6][80] = 16'h0000;
	mel_filter_coefs[6][81] = 16'h0000;
	mel_filter_coefs[6][82] = 16'h0000;
	mel_filter_coefs[6][83] = 16'h0000;
	mel_filter_coefs[6][84] = 16'h0000;
	mel_filter_coefs[6][85] = 16'h0000;
	mel_filter_coefs[6][86] = 16'h0000;
	mel_filter_coefs[6][87] = 16'h0000;
	mel_filter_coefs[6][88] = 16'h0000;
	mel_filter_coefs[6][89] = 16'h0000;
	mel_filter_coefs[6][90] = 16'h0000;
	mel_filter_coefs[6][91] = 16'h0000;
	mel_filter_coefs[6][92] = 16'h0000;
	mel_filter_coefs[6][93] = 16'h0000;
	mel_filter_coefs[6][94] = 16'h0000;
	mel_filter_coefs[6][95] = 16'h0000;
	mel_filter_coefs[6][96] = 16'h0000;
	mel_filter_coefs[6][97] = 16'h0000;
	mel_filter_coefs[6][98] = 16'h0000;
	mel_filter_coefs[6][99] = 16'h0000;
	mel_filter_coefs[6][100] = 16'h0000;
	mel_filter_coefs[6][101] = 16'h0000;
	mel_filter_coefs[6][102] = 16'h0000;
	mel_filter_coefs[6][103] = 16'h0000;
	mel_filter_coefs[6][104] = 16'h0000;
	mel_filter_coefs[6][105] = 16'h0000;
	mel_filter_coefs[6][106] = 16'h0000;
	mel_filter_coefs[6][107] = 16'h0000;
	mel_filter_coefs[6][108] = 16'h0000;
	mel_filter_coefs[6][109] = 16'h0000;
	mel_filter_coefs[6][110] = 16'h0000;
	mel_filter_coefs[6][111] = 16'h0000;
	mel_filter_coefs[6][112] = 16'h0000;
	mel_filter_coefs[6][113] = 16'h0000;
	mel_filter_coefs[6][114] = 16'h0000;
	mel_filter_coefs[6][115] = 16'h0000;
	mel_filter_coefs[6][116] = 16'h0000;
	mel_filter_coefs[6][117] = 16'h0000;
	mel_filter_coefs[6][118] = 16'h0000;
	mel_filter_coefs[6][119] = 16'h0000;
	mel_filter_coefs[6][120] = 16'h0000;
	mel_filter_coefs[6][121] = 16'h0000;
	mel_filter_coefs[6][122] = 16'h0000;
	mel_filter_coefs[6][123] = 16'h0000;
	mel_filter_coefs[6][124] = 16'h0000;
	mel_filter_coefs[6][125] = 16'h0000;
	mel_filter_coefs[6][126] = 16'h0000;
	mel_filter_coefs[6][127] = 16'h0000;
	mel_filter_coefs[6][128] = 16'h0000;
	mel_filter_coefs[6][129] = 16'h0000;
	mel_filter_coefs[6][130] = 16'h0000;
	mel_filter_coefs[6][131] = 16'h0000;
	mel_filter_coefs[6][132] = 16'h0000;
	mel_filter_coefs[6][133] = 16'h0000;
	mel_filter_coefs[6][134] = 16'h0000;
	mel_filter_coefs[6][135] = 16'h0000;
	mel_filter_coefs[6][136] = 16'h0000;
	mel_filter_coefs[6][137] = 16'h0000;
	mel_filter_coefs[6][138] = 16'h0000;
	mel_filter_coefs[6][139] = 16'h0000;
	mel_filter_coefs[6][140] = 16'h0000;
	mel_filter_coefs[6][141] = 16'h0000;
	mel_filter_coefs[6][142] = 16'h0000;
	mel_filter_coefs[6][143] = 16'h0000;
	mel_filter_coefs[6][144] = 16'h0000;
	mel_filter_coefs[6][145] = 16'h0000;
	mel_filter_coefs[6][146] = 16'h0000;
	mel_filter_coefs[6][147] = 16'h0000;
	mel_filter_coefs[6][148] = 16'h0000;
	mel_filter_coefs[6][149] = 16'h0000;
	mel_filter_coefs[6][150] = 16'h0000;
	mel_filter_coefs[6][151] = 16'h0000;
	mel_filter_coefs[6][152] = 16'h0000;
	mel_filter_coefs[6][153] = 16'h0000;
	mel_filter_coefs[6][154] = 16'h0000;
	mel_filter_coefs[6][155] = 16'h0000;
	mel_filter_coefs[6][156] = 16'h0000;
	mel_filter_coefs[6][157] = 16'h0000;
	mel_filter_coefs[6][158] = 16'h0000;
	mel_filter_coefs[6][159] = 16'h0000;
	mel_filter_coefs[6][160] = 16'h0000;
	mel_filter_coefs[6][161] = 16'h0000;
	mel_filter_coefs[6][162] = 16'h0000;
	mel_filter_coefs[6][163] = 16'h0000;
	mel_filter_coefs[6][164] = 16'h0000;
	mel_filter_coefs[6][165] = 16'h0000;
	mel_filter_coefs[6][166] = 16'h0000;
	mel_filter_coefs[6][167] = 16'h0000;
	mel_filter_coefs[6][168] = 16'h0000;
	mel_filter_coefs[6][169] = 16'h0000;
	mel_filter_coefs[6][170] = 16'h0000;
	mel_filter_coefs[6][171] = 16'h0000;
	mel_filter_coefs[6][172] = 16'h0000;
	mel_filter_coefs[6][173] = 16'h0000;
	mel_filter_coefs[6][174] = 16'h0000;
	mel_filter_coefs[6][175] = 16'h0000;
	mel_filter_coefs[6][176] = 16'h0000;
	mel_filter_coefs[6][177] = 16'h0000;
	mel_filter_coefs[6][178] = 16'h0000;
	mel_filter_coefs[6][179] = 16'h0000;
	mel_filter_coefs[6][180] = 16'h0000;
	mel_filter_coefs[6][181] = 16'h0000;
	mel_filter_coefs[6][182] = 16'h0000;
	mel_filter_coefs[6][183] = 16'h0000;
	mel_filter_coefs[6][184] = 16'h0000;
	mel_filter_coefs[6][185] = 16'h0000;
	mel_filter_coefs[6][186] = 16'h0000;
	mel_filter_coefs[6][187] = 16'h0000;
	mel_filter_coefs[6][188] = 16'h0000;
	mel_filter_coefs[6][189] = 16'h0000;
	mel_filter_coefs[6][190] = 16'h0000;
	mel_filter_coefs[6][191] = 16'h0000;
	mel_filter_coefs[6][192] = 16'h0000;
	mel_filter_coefs[6][193] = 16'h0000;
	mel_filter_coefs[6][194] = 16'h0000;
	mel_filter_coefs[6][195] = 16'h0000;
	mel_filter_coefs[6][196] = 16'h0000;
	mel_filter_coefs[6][197] = 16'h0000;
	mel_filter_coefs[6][198] = 16'h0000;
	mel_filter_coefs[6][199] = 16'h0000;
	mel_filter_coefs[6][200] = 16'h0000;
	mel_filter_coefs[6][201] = 16'h0000;
	mel_filter_coefs[6][202] = 16'h0000;
	mel_filter_coefs[6][203] = 16'h0000;
	mel_filter_coefs[6][204] = 16'h0000;
	mel_filter_coefs[6][205] = 16'h0000;
	mel_filter_coefs[6][206] = 16'h0000;
	mel_filter_coefs[6][207] = 16'h0000;
	mel_filter_coefs[6][208] = 16'h0000;
	mel_filter_coefs[6][209] = 16'h0000;
	mel_filter_coefs[6][210] = 16'h0000;
	mel_filter_coefs[6][211] = 16'h0000;
	mel_filter_coefs[6][212] = 16'h0000;
	mel_filter_coefs[6][213] = 16'h0000;
	mel_filter_coefs[6][214] = 16'h0000;
	mel_filter_coefs[6][215] = 16'h0000;
	mel_filter_coefs[6][216] = 16'h0000;
	mel_filter_coefs[6][217] = 16'h0000;
	mel_filter_coefs[6][218] = 16'h0000;
	mel_filter_coefs[6][219] = 16'h0000;
	mel_filter_coefs[6][220] = 16'h0000;
	mel_filter_coefs[6][221] = 16'h0000;
	mel_filter_coefs[6][222] = 16'h0000;
	mel_filter_coefs[6][223] = 16'h0000;
	mel_filter_coefs[6][224] = 16'h0000;
	mel_filter_coefs[6][225] = 16'h0000;
	mel_filter_coefs[6][226] = 16'h0000;
	mel_filter_coefs[6][227] = 16'h0000;
	mel_filter_coefs[6][228] = 16'h0000;
	mel_filter_coefs[6][229] = 16'h0000;
	mel_filter_coefs[6][230] = 16'h0000;
	mel_filter_coefs[6][231] = 16'h0000;
	mel_filter_coefs[6][232] = 16'h0000;
	mel_filter_coefs[6][233] = 16'h0000;
	mel_filter_coefs[6][234] = 16'h0000;
	mel_filter_coefs[6][235] = 16'h0000;
	mel_filter_coefs[6][236] = 16'h0000;
	mel_filter_coefs[6][237] = 16'h0000;
	mel_filter_coefs[6][238] = 16'h0000;
	mel_filter_coefs[6][239] = 16'h0000;
	mel_filter_coefs[6][240] = 16'h0000;
	mel_filter_coefs[6][241] = 16'h0000;
	mel_filter_coefs[6][242] = 16'h0000;
	mel_filter_coefs[6][243] = 16'h0000;
	mel_filter_coefs[6][244] = 16'h0000;
	mel_filter_coefs[6][245] = 16'h0000;
	mel_filter_coefs[6][246] = 16'h0000;
	mel_filter_coefs[6][247] = 16'h0000;
	mel_filter_coefs[6][248] = 16'h0000;
	mel_filter_coefs[6][249] = 16'h0000;
	mel_filter_coefs[6][250] = 16'h0000;
	mel_filter_coefs[6][251] = 16'h0000;
	mel_filter_coefs[6][252] = 16'h0000;
	mel_filter_coefs[6][253] = 16'h0000;
	mel_filter_coefs[6][254] = 16'h0000;
	mel_filter_coefs[6][255] = 16'h0000;
	mel_filter_coefs[7][0] = 16'h0000;
	mel_filter_coefs[7][1] = 16'h0000;
	mel_filter_coefs[7][2] = 16'h0000;
	mel_filter_coefs[7][3] = 16'h0000;
	mel_filter_coefs[7][4] = 16'h0000;
	mel_filter_coefs[7][5] = 16'h0000;
	mel_filter_coefs[7][6] = 16'h0000;
	mel_filter_coefs[7][7] = 16'h0000;
	mel_filter_coefs[7][8] = 16'h0000;
	mel_filter_coefs[7][9] = 16'h0000;
	mel_filter_coefs[7][10] = 16'h0000;
	mel_filter_coefs[7][11] = 16'h0000;
	mel_filter_coefs[7][12] = 16'h003E;
	mel_filter_coefs[7][13] = 16'h3B18;
	mel_filter_coefs[7][14] = 16'h75F3;
	mel_filter_coefs[7][15] = 16'h521B;
	mel_filter_coefs[7][16] = 16'h1AC3;
	mel_filter_coefs[7][17] = 16'h0000;
	mel_filter_coefs[7][18] = 16'h0000;
	mel_filter_coefs[7][19] = 16'h0000;
	mel_filter_coefs[7][20] = 16'h0000;
	mel_filter_coefs[7][21] = 16'h0000;
	mel_filter_coefs[7][22] = 16'h0000;
	mel_filter_coefs[7][23] = 16'h0000;
	mel_filter_coefs[7][24] = 16'h0000;
	mel_filter_coefs[7][25] = 16'h0000;
	mel_filter_coefs[7][26] = 16'h0000;
	mel_filter_coefs[7][27] = 16'h0000;
	mel_filter_coefs[7][28] = 16'h0000;
	mel_filter_coefs[7][29] = 16'h0000;
	mel_filter_coefs[7][30] = 16'h0000;
	mel_filter_coefs[7][31] = 16'h0000;
	mel_filter_coefs[7][32] = 16'h0000;
	mel_filter_coefs[7][33] = 16'h0000;
	mel_filter_coefs[7][34] = 16'h0000;
	mel_filter_coefs[7][35] = 16'h0000;
	mel_filter_coefs[7][36] = 16'h0000;
	mel_filter_coefs[7][37] = 16'h0000;
	mel_filter_coefs[7][38] = 16'h0000;
	mel_filter_coefs[7][39] = 16'h0000;
	mel_filter_coefs[7][40] = 16'h0000;
	mel_filter_coefs[7][41] = 16'h0000;
	mel_filter_coefs[7][42] = 16'h0000;
	mel_filter_coefs[7][43] = 16'h0000;
	mel_filter_coefs[7][44] = 16'h0000;
	mel_filter_coefs[7][45] = 16'h0000;
	mel_filter_coefs[7][46] = 16'h0000;
	mel_filter_coefs[7][47] = 16'h0000;
	mel_filter_coefs[7][48] = 16'h0000;
	mel_filter_coefs[7][49] = 16'h0000;
	mel_filter_coefs[7][50] = 16'h0000;
	mel_filter_coefs[7][51] = 16'h0000;
	mel_filter_coefs[7][52] = 16'h0000;
	mel_filter_coefs[7][53] = 16'h0000;
	mel_filter_coefs[7][54] = 16'h0000;
	mel_filter_coefs[7][55] = 16'h0000;
	mel_filter_coefs[7][56] = 16'h0000;
	mel_filter_coefs[7][57] = 16'h0000;
	mel_filter_coefs[7][58] = 16'h0000;
	mel_filter_coefs[7][59] = 16'h0000;
	mel_filter_coefs[7][60] = 16'h0000;
	mel_filter_coefs[7][61] = 16'h0000;
	mel_filter_coefs[7][62] = 16'h0000;
	mel_filter_coefs[7][63] = 16'h0000;
	mel_filter_coefs[7][64] = 16'h0000;
	mel_filter_coefs[7][65] = 16'h0000;
	mel_filter_coefs[7][66] = 16'h0000;
	mel_filter_coefs[7][67] = 16'h0000;
	mel_filter_coefs[7][68] = 16'h0000;
	mel_filter_coefs[7][69] = 16'h0000;
	mel_filter_coefs[7][70] = 16'h0000;
	mel_filter_coefs[7][71] = 16'h0000;
	mel_filter_coefs[7][72] = 16'h0000;
	mel_filter_coefs[7][73] = 16'h0000;
	mel_filter_coefs[7][74] = 16'h0000;
	mel_filter_coefs[7][75] = 16'h0000;
	mel_filter_coefs[7][76] = 16'h0000;
	mel_filter_coefs[7][77] = 16'h0000;
	mel_filter_coefs[7][78] = 16'h0000;
	mel_filter_coefs[7][79] = 16'h0000;
	mel_filter_coefs[7][80] = 16'h0000;
	mel_filter_coefs[7][81] = 16'h0000;
	mel_filter_coefs[7][82] = 16'h0000;
	mel_filter_coefs[7][83] = 16'h0000;
	mel_filter_coefs[7][84] = 16'h0000;
	mel_filter_coefs[7][85] = 16'h0000;
	mel_filter_coefs[7][86] = 16'h0000;
	mel_filter_coefs[7][87] = 16'h0000;
	mel_filter_coefs[7][88] = 16'h0000;
	mel_filter_coefs[7][89] = 16'h0000;
	mel_filter_coefs[7][90] = 16'h0000;
	mel_filter_coefs[7][91] = 16'h0000;
	mel_filter_coefs[7][92] = 16'h0000;
	mel_filter_coefs[7][93] = 16'h0000;
	mel_filter_coefs[7][94] = 16'h0000;
	mel_filter_coefs[7][95] = 16'h0000;
	mel_filter_coefs[7][96] = 16'h0000;
	mel_filter_coefs[7][97] = 16'h0000;
	mel_filter_coefs[7][98] = 16'h0000;
	mel_filter_coefs[7][99] = 16'h0000;
	mel_filter_coefs[7][100] = 16'h0000;
	mel_filter_coefs[7][101] = 16'h0000;
	mel_filter_coefs[7][102] = 16'h0000;
	mel_filter_coefs[7][103] = 16'h0000;
	mel_filter_coefs[7][104] = 16'h0000;
	mel_filter_coefs[7][105] = 16'h0000;
	mel_filter_coefs[7][106] = 16'h0000;
	mel_filter_coefs[7][107] = 16'h0000;
	mel_filter_coefs[7][108] = 16'h0000;
	mel_filter_coefs[7][109] = 16'h0000;
	mel_filter_coefs[7][110] = 16'h0000;
	mel_filter_coefs[7][111] = 16'h0000;
	mel_filter_coefs[7][112] = 16'h0000;
	mel_filter_coefs[7][113] = 16'h0000;
	mel_filter_coefs[7][114] = 16'h0000;
	mel_filter_coefs[7][115] = 16'h0000;
	mel_filter_coefs[7][116] = 16'h0000;
	mel_filter_coefs[7][117] = 16'h0000;
	mel_filter_coefs[7][118] = 16'h0000;
	mel_filter_coefs[7][119] = 16'h0000;
	mel_filter_coefs[7][120] = 16'h0000;
	mel_filter_coefs[7][121] = 16'h0000;
	mel_filter_coefs[7][122] = 16'h0000;
	mel_filter_coefs[7][123] = 16'h0000;
	mel_filter_coefs[7][124] = 16'h0000;
	mel_filter_coefs[7][125] = 16'h0000;
	mel_filter_coefs[7][126] = 16'h0000;
	mel_filter_coefs[7][127] = 16'h0000;
	mel_filter_coefs[7][128] = 16'h0000;
	mel_filter_coefs[7][129] = 16'h0000;
	mel_filter_coefs[7][130] = 16'h0000;
	mel_filter_coefs[7][131] = 16'h0000;
	mel_filter_coefs[7][132] = 16'h0000;
	mel_filter_coefs[7][133] = 16'h0000;
	mel_filter_coefs[7][134] = 16'h0000;
	mel_filter_coefs[7][135] = 16'h0000;
	mel_filter_coefs[7][136] = 16'h0000;
	mel_filter_coefs[7][137] = 16'h0000;
	mel_filter_coefs[7][138] = 16'h0000;
	mel_filter_coefs[7][139] = 16'h0000;
	mel_filter_coefs[7][140] = 16'h0000;
	mel_filter_coefs[7][141] = 16'h0000;
	mel_filter_coefs[7][142] = 16'h0000;
	mel_filter_coefs[7][143] = 16'h0000;
	mel_filter_coefs[7][144] = 16'h0000;
	mel_filter_coefs[7][145] = 16'h0000;
	mel_filter_coefs[7][146] = 16'h0000;
	mel_filter_coefs[7][147] = 16'h0000;
	mel_filter_coefs[7][148] = 16'h0000;
	mel_filter_coefs[7][149] = 16'h0000;
	mel_filter_coefs[7][150] = 16'h0000;
	mel_filter_coefs[7][151] = 16'h0000;
	mel_filter_coefs[7][152] = 16'h0000;
	mel_filter_coefs[7][153] = 16'h0000;
	mel_filter_coefs[7][154] = 16'h0000;
	mel_filter_coefs[7][155] = 16'h0000;
	mel_filter_coefs[7][156] = 16'h0000;
	mel_filter_coefs[7][157] = 16'h0000;
	mel_filter_coefs[7][158] = 16'h0000;
	mel_filter_coefs[7][159] = 16'h0000;
	mel_filter_coefs[7][160] = 16'h0000;
	mel_filter_coefs[7][161] = 16'h0000;
	mel_filter_coefs[7][162] = 16'h0000;
	mel_filter_coefs[7][163] = 16'h0000;
	mel_filter_coefs[7][164] = 16'h0000;
	mel_filter_coefs[7][165] = 16'h0000;
	mel_filter_coefs[7][166] = 16'h0000;
	mel_filter_coefs[7][167] = 16'h0000;
	mel_filter_coefs[7][168] = 16'h0000;
	mel_filter_coefs[7][169] = 16'h0000;
	mel_filter_coefs[7][170] = 16'h0000;
	mel_filter_coefs[7][171] = 16'h0000;
	mel_filter_coefs[7][172] = 16'h0000;
	mel_filter_coefs[7][173] = 16'h0000;
	mel_filter_coefs[7][174] = 16'h0000;
	mel_filter_coefs[7][175] = 16'h0000;
	mel_filter_coefs[7][176] = 16'h0000;
	mel_filter_coefs[7][177] = 16'h0000;
	mel_filter_coefs[7][178] = 16'h0000;
	mel_filter_coefs[7][179] = 16'h0000;
	mel_filter_coefs[7][180] = 16'h0000;
	mel_filter_coefs[7][181] = 16'h0000;
	mel_filter_coefs[7][182] = 16'h0000;
	mel_filter_coefs[7][183] = 16'h0000;
	mel_filter_coefs[7][184] = 16'h0000;
	mel_filter_coefs[7][185] = 16'h0000;
	mel_filter_coefs[7][186] = 16'h0000;
	mel_filter_coefs[7][187] = 16'h0000;
	mel_filter_coefs[7][188] = 16'h0000;
	mel_filter_coefs[7][189] = 16'h0000;
	mel_filter_coefs[7][190] = 16'h0000;
	mel_filter_coefs[7][191] = 16'h0000;
	mel_filter_coefs[7][192] = 16'h0000;
	mel_filter_coefs[7][193] = 16'h0000;
	mel_filter_coefs[7][194] = 16'h0000;
	mel_filter_coefs[7][195] = 16'h0000;
	mel_filter_coefs[7][196] = 16'h0000;
	mel_filter_coefs[7][197] = 16'h0000;
	mel_filter_coefs[7][198] = 16'h0000;
	mel_filter_coefs[7][199] = 16'h0000;
	mel_filter_coefs[7][200] = 16'h0000;
	mel_filter_coefs[7][201] = 16'h0000;
	mel_filter_coefs[7][202] = 16'h0000;
	mel_filter_coefs[7][203] = 16'h0000;
	mel_filter_coefs[7][204] = 16'h0000;
	mel_filter_coefs[7][205] = 16'h0000;
	mel_filter_coefs[7][206] = 16'h0000;
	mel_filter_coefs[7][207] = 16'h0000;
	mel_filter_coefs[7][208] = 16'h0000;
	mel_filter_coefs[7][209] = 16'h0000;
	mel_filter_coefs[7][210] = 16'h0000;
	mel_filter_coefs[7][211] = 16'h0000;
	mel_filter_coefs[7][212] = 16'h0000;
	mel_filter_coefs[7][213] = 16'h0000;
	mel_filter_coefs[7][214] = 16'h0000;
	mel_filter_coefs[7][215] = 16'h0000;
	mel_filter_coefs[7][216] = 16'h0000;
	mel_filter_coefs[7][217] = 16'h0000;
	mel_filter_coefs[7][218] = 16'h0000;
	mel_filter_coefs[7][219] = 16'h0000;
	mel_filter_coefs[7][220] = 16'h0000;
	mel_filter_coefs[7][221] = 16'h0000;
	mel_filter_coefs[7][222] = 16'h0000;
	mel_filter_coefs[7][223] = 16'h0000;
	mel_filter_coefs[7][224] = 16'h0000;
	mel_filter_coefs[7][225] = 16'h0000;
	mel_filter_coefs[7][226] = 16'h0000;
	mel_filter_coefs[7][227] = 16'h0000;
	mel_filter_coefs[7][228] = 16'h0000;
	mel_filter_coefs[7][229] = 16'h0000;
	mel_filter_coefs[7][230] = 16'h0000;
	mel_filter_coefs[7][231] = 16'h0000;
	mel_filter_coefs[7][232] = 16'h0000;
	mel_filter_coefs[7][233] = 16'h0000;
	mel_filter_coefs[7][234] = 16'h0000;
	mel_filter_coefs[7][235] = 16'h0000;
	mel_filter_coefs[7][236] = 16'h0000;
	mel_filter_coefs[7][237] = 16'h0000;
	mel_filter_coefs[7][238] = 16'h0000;
	mel_filter_coefs[7][239] = 16'h0000;
	mel_filter_coefs[7][240] = 16'h0000;
	mel_filter_coefs[7][241] = 16'h0000;
	mel_filter_coefs[7][242] = 16'h0000;
	mel_filter_coefs[7][243] = 16'h0000;
	mel_filter_coefs[7][244] = 16'h0000;
	mel_filter_coefs[7][245] = 16'h0000;
	mel_filter_coefs[7][246] = 16'h0000;
	mel_filter_coefs[7][247] = 16'h0000;
	mel_filter_coefs[7][248] = 16'h0000;
	mel_filter_coefs[7][249] = 16'h0000;
	mel_filter_coefs[7][250] = 16'h0000;
	mel_filter_coefs[7][251] = 16'h0000;
	mel_filter_coefs[7][252] = 16'h0000;
	mel_filter_coefs[7][253] = 16'h0000;
	mel_filter_coefs[7][254] = 16'h0000;
	mel_filter_coefs[7][255] = 16'h0000;
	mel_filter_coefs[8][0] = 16'h0000;
	mel_filter_coefs[8][1] = 16'h0000;
	mel_filter_coefs[8][2] = 16'h0000;
	mel_filter_coefs[8][3] = 16'h0000;
	mel_filter_coefs[8][4] = 16'h0000;
	mel_filter_coefs[8][5] = 16'h0000;
	mel_filter_coefs[8][6] = 16'h0000;
	mel_filter_coefs[8][7] = 16'h0000;
	mel_filter_coefs[8][8] = 16'h0000;
	mel_filter_coefs[8][9] = 16'h0000;
	mel_filter_coefs[8][10] = 16'h0000;
	mel_filter_coefs[8][11] = 16'h0000;
	mel_filter_coefs[8][12] = 16'h0000;
	mel_filter_coefs[8][13] = 16'h0000;
	mel_filter_coefs[8][14] = 16'h0000;
	mel_filter_coefs[8][15] = 16'h2DE5;
	mel_filter_coefs[8][16] = 16'h653D;
	mel_filter_coefs[8][17] = 16'h651E;
	mel_filter_coefs[8][18] = 16'h3112;
	mel_filter_coefs[8][19] = 16'h0000;
	mel_filter_coefs[8][20] = 16'h0000;
	mel_filter_coefs[8][21] = 16'h0000;
	mel_filter_coefs[8][22] = 16'h0000;
	mel_filter_coefs[8][23] = 16'h0000;
	mel_filter_coefs[8][24] = 16'h0000;
	mel_filter_coefs[8][25] = 16'h0000;
	mel_filter_coefs[8][26] = 16'h0000;
	mel_filter_coefs[8][27] = 16'h0000;
	mel_filter_coefs[8][28] = 16'h0000;
	mel_filter_coefs[8][29] = 16'h0000;
	mel_filter_coefs[8][30] = 16'h0000;
	mel_filter_coefs[8][31] = 16'h0000;
	mel_filter_coefs[8][32] = 16'h0000;
	mel_filter_coefs[8][33] = 16'h0000;
	mel_filter_coefs[8][34] = 16'h0000;
	mel_filter_coefs[8][35] = 16'h0000;
	mel_filter_coefs[8][36] = 16'h0000;
	mel_filter_coefs[8][37] = 16'h0000;
	mel_filter_coefs[8][38] = 16'h0000;
	mel_filter_coefs[8][39] = 16'h0000;
	mel_filter_coefs[8][40] = 16'h0000;
	mel_filter_coefs[8][41] = 16'h0000;
	mel_filter_coefs[8][42] = 16'h0000;
	mel_filter_coefs[8][43] = 16'h0000;
	mel_filter_coefs[8][44] = 16'h0000;
	mel_filter_coefs[8][45] = 16'h0000;
	mel_filter_coefs[8][46] = 16'h0000;
	mel_filter_coefs[8][47] = 16'h0000;
	mel_filter_coefs[8][48] = 16'h0000;
	mel_filter_coefs[8][49] = 16'h0000;
	mel_filter_coefs[8][50] = 16'h0000;
	mel_filter_coefs[8][51] = 16'h0000;
	mel_filter_coefs[8][52] = 16'h0000;
	mel_filter_coefs[8][53] = 16'h0000;
	mel_filter_coefs[8][54] = 16'h0000;
	mel_filter_coefs[8][55] = 16'h0000;
	mel_filter_coefs[8][56] = 16'h0000;
	mel_filter_coefs[8][57] = 16'h0000;
	mel_filter_coefs[8][58] = 16'h0000;
	mel_filter_coefs[8][59] = 16'h0000;
	mel_filter_coefs[8][60] = 16'h0000;
	mel_filter_coefs[8][61] = 16'h0000;
	mel_filter_coefs[8][62] = 16'h0000;
	mel_filter_coefs[8][63] = 16'h0000;
	mel_filter_coefs[8][64] = 16'h0000;
	mel_filter_coefs[8][65] = 16'h0000;
	mel_filter_coefs[8][66] = 16'h0000;
	mel_filter_coefs[8][67] = 16'h0000;
	mel_filter_coefs[8][68] = 16'h0000;
	mel_filter_coefs[8][69] = 16'h0000;
	mel_filter_coefs[8][70] = 16'h0000;
	mel_filter_coefs[8][71] = 16'h0000;
	mel_filter_coefs[8][72] = 16'h0000;
	mel_filter_coefs[8][73] = 16'h0000;
	mel_filter_coefs[8][74] = 16'h0000;
	mel_filter_coefs[8][75] = 16'h0000;
	mel_filter_coefs[8][76] = 16'h0000;
	mel_filter_coefs[8][77] = 16'h0000;
	mel_filter_coefs[8][78] = 16'h0000;
	mel_filter_coefs[8][79] = 16'h0000;
	mel_filter_coefs[8][80] = 16'h0000;
	mel_filter_coefs[8][81] = 16'h0000;
	mel_filter_coefs[8][82] = 16'h0000;
	mel_filter_coefs[8][83] = 16'h0000;
	mel_filter_coefs[8][84] = 16'h0000;
	mel_filter_coefs[8][85] = 16'h0000;
	mel_filter_coefs[8][86] = 16'h0000;
	mel_filter_coefs[8][87] = 16'h0000;
	mel_filter_coefs[8][88] = 16'h0000;
	mel_filter_coefs[8][89] = 16'h0000;
	mel_filter_coefs[8][90] = 16'h0000;
	mel_filter_coefs[8][91] = 16'h0000;
	mel_filter_coefs[8][92] = 16'h0000;
	mel_filter_coefs[8][93] = 16'h0000;
	mel_filter_coefs[8][94] = 16'h0000;
	mel_filter_coefs[8][95] = 16'h0000;
	mel_filter_coefs[8][96] = 16'h0000;
	mel_filter_coefs[8][97] = 16'h0000;
	mel_filter_coefs[8][98] = 16'h0000;
	mel_filter_coefs[8][99] = 16'h0000;
	mel_filter_coefs[8][100] = 16'h0000;
	mel_filter_coefs[8][101] = 16'h0000;
	mel_filter_coefs[8][102] = 16'h0000;
	mel_filter_coefs[8][103] = 16'h0000;
	mel_filter_coefs[8][104] = 16'h0000;
	mel_filter_coefs[8][105] = 16'h0000;
	mel_filter_coefs[8][106] = 16'h0000;
	mel_filter_coefs[8][107] = 16'h0000;
	mel_filter_coefs[8][108] = 16'h0000;
	mel_filter_coefs[8][109] = 16'h0000;
	mel_filter_coefs[8][110] = 16'h0000;
	mel_filter_coefs[8][111] = 16'h0000;
	mel_filter_coefs[8][112] = 16'h0000;
	mel_filter_coefs[8][113] = 16'h0000;
	mel_filter_coefs[8][114] = 16'h0000;
	mel_filter_coefs[8][115] = 16'h0000;
	mel_filter_coefs[8][116] = 16'h0000;
	mel_filter_coefs[8][117] = 16'h0000;
	mel_filter_coefs[8][118] = 16'h0000;
	mel_filter_coefs[8][119] = 16'h0000;
	mel_filter_coefs[8][120] = 16'h0000;
	mel_filter_coefs[8][121] = 16'h0000;
	mel_filter_coefs[8][122] = 16'h0000;
	mel_filter_coefs[8][123] = 16'h0000;
	mel_filter_coefs[8][124] = 16'h0000;
	mel_filter_coefs[8][125] = 16'h0000;
	mel_filter_coefs[8][126] = 16'h0000;
	mel_filter_coefs[8][127] = 16'h0000;
	mel_filter_coefs[8][128] = 16'h0000;
	mel_filter_coefs[8][129] = 16'h0000;
	mel_filter_coefs[8][130] = 16'h0000;
	mel_filter_coefs[8][131] = 16'h0000;
	mel_filter_coefs[8][132] = 16'h0000;
	mel_filter_coefs[8][133] = 16'h0000;
	mel_filter_coefs[8][134] = 16'h0000;
	mel_filter_coefs[8][135] = 16'h0000;
	mel_filter_coefs[8][136] = 16'h0000;
	mel_filter_coefs[8][137] = 16'h0000;
	mel_filter_coefs[8][138] = 16'h0000;
	mel_filter_coefs[8][139] = 16'h0000;
	mel_filter_coefs[8][140] = 16'h0000;
	mel_filter_coefs[8][141] = 16'h0000;
	mel_filter_coefs[8][142] = 16'h0000;
	mel_filter_coefs[8][143] = 16'h0000;
	mel_filter_coefs[8][144] = 16'h0000;
	mel_filter_coefs[8][145] = 16'h0000;
	mel_filter_coefs[8][146] = 16'h0000;
	mel_filter_coefs[8][147] = 16'h0000;
	mel_filter_coefs[8][148] = 16'h0000;
	mel_filter_coefs[8][149] = 16'h0000;
	mel_filter_coefs[8][150] = 16'h0000;
	mel_filter_coefs[8][151] = 16'h0000;
	mel_filter_coefs[8][152] = 16'h0000;
	mel_filter_coefs[8][153] = 16'h0000;
	mel_filter_coefs[8][154] = 16'h0000;
	mel_filter_coefs[8][155] = 16'h0000;
	mel_filter_coefs[8][156] = 16'h0000;
	mel_filter_coefs[8][157] = 16'h0000;
	mel_filter_coefs[8][158] = 16'h0000;
	mel_filter_coefs[8][159] = 16'h0000;
	mel_filter_coefs[8][160] = 16'h0000;
	mel_filter_coefs[8][161] = 16'h0000;
	mel_filter_coefs[8][162] = 16'h0000;
	mel_filter_coefs[8][163] = 16'h0000;
	mel_filter_coefs[8][164] = 16'h0000;
	mel_filter_coefs[8][165] = 16'h0000;
	mel_filter_coefs[8][166] = 16'h0000;
	mel_filter_coefs[8][167] = 16'h0000;
	mel_filter_coefs[8][168] = 16'h0000;
	mel_filter_coefs[8][169] = 16'h0000;
	mel_filter_coefs[8][170] = 16'h0000;
	mel_filter_coefs[8][171] = 16'h0000;
	mel_filter_coefs[8][172] = 16'h0000;
	mel_filter_coefs[8][173] = 16'h0000;
	mel_filter_coefs[8][174] = 16'h0000;
	mel_filter_coefs[8][175] = 16'h0000;
	mel_filter_coefs[8][176] = 16'h0000;
	mel_filter_coefs[8][177] = 16'h0000;
	mel_filter_coefs[8][178] = 16'h0000;
	mel_filter_coefs[8][179] = 16'h0000;
	mel_filter_coefs[8][180] = 16'h0000;
	mel_filter_coefs[8][181] = 16'h0000;
	mel_filter_coefs[8][182] = 16'h0000;
	mel_filter_coefs[8][183] = 16'h0000;
	mel_filter_coefs[8][184] = 16'h0000;
	mel_filter_coefs[8][185] = 16'h0000;
	mel_filter_coefs[8][186] = 16'h0000;
	mel_filter_coefs[8][187] = 16'h0000;
	mel_filter_coefs[8][188] = 16'h0000;
	mel_filter_coefs[8][189] = 16'h0000;
	mel_filter_coefs[8][190] = 16'h0000;
	mel_filter_coefs[8][191] = 16'h0000;
	mel_filter_coefs[8][192] = 16'h0000;
	mel_filter_coefs[8][193] = 16'h0000;
	mel_filter_coefs[8][194] = 16'h0000;
	mel_filter_coefs[8][195] = 16'h0000;
	mel_filter_coefs[8][196] = 16'h0000;
	mel_filter_coefs[8][197] = 16'h0000;
	mel_filter_coefs[8][198] = 16'h0000;
	mel_filter_coefs[8][199] = 16'h0000;
	mel_filter_coefs[8][200] = 16'h0000;
	mel_filter_coefs[8][201] = 16'h0000;
	mel_filter_coefs[8][202] = 16'h0000;
	mel_filter_coefs[8][203] = 16'h0000;
	mel_filter_coefs[8][204] = 16'h0000;
	mel_filter_coefs[8][205] = 16'h0000;
	mel_filter_coefs[8][206] = 16'h0000;
	mel_filter_coefs[8][207] = 16'h0000;
	mel_filter_coefs[8][208] = 16'h0000;
	mel_filter_coefs[8][209] = 16'h0000;
	mel_filter_coefs[8][210] = 16'h0000;
	mel_filter_coefs[8][211] = 16'h0000;
	mel_filter_coefs[8][212] = 16'h0000;
	mel_filter_coefs[8][213] = 16'h0000;
	mel_filter_coefs[8][214] = 16'h0000;
	mel_filter_coefs[8][215] = 16'h0000;
	mel_filter_coefs[8][216] = 16'h0000;
	mel_filter_coefs[8][217] = 16'h0000;
	mel_filter_coefs[8][218] = 16'h0000;
	mel_filter_coefs[8][219] = 16'h0000;
	mel_filter_coefs[8][220] = 16'h0000;
	mel_filter_coefs[8][221] = 16'h0000;
	mel_filter_coefs[8][222] = 16'h0000;
	mel_filter_coefs[8][223] = 16'h0000;
	mel_filter_coefs[8][224] = 16'h0000;
	mel_filter_coefs[8][225] = 16'h0000;
	mel_filter_coefs[8][226] = 16'h0000;
	mel_filter_coefs[8][227] = 16'h0000;
	mel_filter_coefs[8][228] = 16'h0000;
	mel_filter_coefs[8][229] = 16'h0000;
	mel_filter_coefs[8][230] = 16'h0000;
	mel_filter_coefs[8][231] = 16'h0000;
	mel_filter_coefs[8][232] = 16'h0000;
	mel_filter_coefs[8][233] = 16'h0000;
	mel_filter_coefs[8][234] = 16'h0000;
	mel_filter_coefs[8][235] = 16'h0000;
	mel_filter_coefs[8][236] = 16'h0000;
	mel_filter_coefs[8][237] = 16'h0000;
	mel_filter_coefs[8][238] = 16'h0000;
	mel_filter_coefs[8][239] = 16'h0000;
	mel_filter_coefs[8][240] = 16'h0000;
	mel_filter_coefs[8][241] = 16'h0000;
	mel_filter_coefs[8][242] = 16'h0000;
	mel_filter_coefs[8][243] = 16'h0000;
	mel_filter_coefs[8][244] = 16'h0000;
	mel_filter_coefs[8][245] = 16'h0000;
	mel_filter_coefs[8][246] = 16'h0000;
	mel_filter_coefs[8][247] = 16'h0000;
	mel_filter_coefs[8][248] = 16'h0000;
	mel_filter_coefs[8][249] = 16'h0000;
	mel_filter_coefs[8][250] = 16'h0000;
	mel_filter_coefs[8][251] = 16'h0000;
	mel_filter_coefs[8][252] = 16'h0000;
	mel_filter_coefs[8][253] = 16'h0000;
	mel_filter_coefs[8][254] = 16'h0000;
	mel_filter_coefs[8][255] = 16'h0000;
	mel_filter_coefs[9][0] = 16'h0000;
	mel_filter_coefs[9][1] = 16'h0000;
	mel_filter_coefs[9][2] = 16'h0000;
	mel_filter_coefs[9][3] = 16'h0000;
	mel_filter_coefs[9][4] = 16'h0000;
	mel_filter_coefs[9][5] = 16'h0000;
	mel_filter_coefs[9][6] = 16'h0000;
	mel_filter_coefs[9][7] = 16'h0000;
	mel_filter_coefs[9][8] = 16'h0000;
	mel_filter_coefs[9][9] = 16'h0000;
	mel_filter_coefs[9][10] = 16'h0000;
	mel_filter_coefs[9][11] = 16'h0000;
	mel_filter_coefs[9][12] = 16'h0000;
	mel_filter_coefs[9][13] = 16'h0000;
	mel_filter_coefs[9][14] = 16'h0000;
	mel_filter_coefs[9][15] = 16'h0000;
	mel_filter_coefs[9][16] = 16'h0000;
	mel_filter_coefs[9][17] = 16'h1AE2;
	mel_filter_coefs[9][18] = 16'h4EEE;
	mel_filter_coefs[9][19] = 16'h7D34;
	mel_filter_coefs[9][20] = 16'h4C42;
	mel_filter_coefs[9][21] = 16'h1B51;
	mel_filter_coefs[9][22] = 16'h0000;
	mel_filter_coefs[9][23] = 16'h0000;
	mel_filter_coefs[9][24] = 16'h0000;
	mel_filter_coefs[9][25] = 16'h0000;
	mel_filter_coefs[9][26] = 16'h0000;
	mel_filter_coefs[9][27] = 16'h0000;
	mel_filter_coefs[9][28] = 16'h0000;
	mel_filter_coefs[9][29] = 16'h0000;
	mel_filter_coefs[9][30] = 16'h0000;
	mel_filter_coefs[9][31] = 16'h0000;
	mel_filter_coefs[9][32] = 16'h0000;
	mel_filter_coefs[9][33] = 16'h0000;
	mel_filter_coefs[9][34] = 16'h0000;
	mel_filter_coefs[9][35] = 16'h0000;
	mel_filter_coefs[9][36] = 16'h0000;
	mel_filter_coefs[9][37] = 16'h0000;
	mel_filter_coefs[9][38] = 16'h0000;
	mel_filter_coefs[9][39] = 16'h0000;
	mel_filter_coefs[9][40] = 16'h0000;
	mel_filter_coefs[9][41] = 16'h0000;
	mel_filter_coefs[9][42] = 16'h0000;
	mel_filter_coefs[9][43] = 16'h0000;
	mel_filter_coefs[9][44] = 16'h0000;
	mel_filter_coefs[9][45] = 16'h0000;
	mel_filter_coefs[9][46] = 16'h0000;
	mel_filter_coefs[9][47] = 16'h0000;
	mel_filter_coefs[9][48] = 16'h0000;
	mel_filter_coefs[9][49] = 16'h0000;
	mel_filter_coefs[9][50] = 16'h0000;
	mel_filter_coefs[9][51] = 16'h0000;
	mel_filter_coefs[9][52] = 16'h0000;
	mel_filter_coefs[9][53] = 16'h0000;
	mel_filter_coefs[9][54] = 16'h0000;
	mel_filter_coefs[9][55] = 16'h0000;
	mel_filter_coefs[9][56] = 16'h0000;
	mel_filter_coefs[9][57] = 16'h0000;
	mel_filter_coefs[9][58] = 16'h0000;
	mel_filter_coefs[9][59] = 16'h0000;
	mel_filter_coefs[9][60] = 16'h0000;
	mel_filter_coefs[9][61] = 16'h0000;
	mel_filter_coefs[9][62] = 16'h0000;
	mel_filter_coefs[9][63] = 16'h0000;
	mel_filter_coefs[9][64] = 16'h0000;
	mel_filter_coefs[9][65] = 16'h0000;
	mel_filter_coefs[9][66] = 16'h0000;
	mel_filter_coefs[9][67] = 16'h0000;
	mel_filter_coefs[9][68] = 16'h0000;
	mel_filter_coefs[9][69] = 16'h0000;
	mel_filter_coefs[9][70] = 16'h0000;
	mel_filter_coefs[9][71] = 16'h0000;
	mel_filter_coefs[9][72] = 16'h0000;
	mel_filter_coefs[9][73] = 16'h0000;
	mel_filter_coefs[9][74] = 16'h0000;
	mel_filter_coefs[9][75] = 16'h0000;
	mel_filter_coefs[9][76] = 16'h0000;
	mel_filter_coefs[9][77] = 16'h0000;
	mel_filter_coefs[9][78] = 16'h0000;
	mel_filter_coefs[9][79] = 16'h0000;
	mel_filter_coefs[9][80] = 16'h0000;
	mel_filter_coefs[9][81] = 16'h0000;
	mel_filter_coefs[9][82] = 16'h0000;
	mel_filter_coefs[9][83] = 16'h0000;
	mel_filter_coefs[9][84] = 16'h0000;
	mel_filter_coefs[9][85] = 16'h0000;
	mel_filter_coefs[9][86] = 16'h0000;
	mel_filter_coefs[9][87] = 16'h0000;
	mel_filter_coefs[9][88] = 16'h0000;
	mel_filter_coefs[9][89] = 16'h0000;
	mel_filter_coefs[9][90] = 16'h0000;
	mel_filter_coefs[9][91] = 16'h0000;
	mel_filter_coefs[9][92] = 16'h0000;
	mel_filter_coefs[9][93] = 16'h0000;
	mel_filter_coefs[9][94] = 16'h0000;
	mel_filter_coefs[9][95] = 16'h0000;
	mel_filter_coefs[9][96] = 16'h0000;
	mel_filter_coefs[9][97] = 16'h0000;
	mel_filter_coefs[9][98] = 16'h0000;
	mel_filter_coefs[9][99] = 16'h0000;
	mel_filter_coefs[9][100] = 16'h0000;
	mel_filter_coefs[9][101] = 16'h0000;
	mel_filter_coefs[9][102] = 16'h0000;
	mel_filter_coefs[9][103] = 16'h0000;
	mel_filter_coefs[9][104] = 16'h0000;
	mel_filter_coefs[9][105] = 16'h0000;
	mel_filter_coefs[9][106] = 16'h0000;
	mel_filter_coefs[9][107] = 16'h0000;
	mel_filter_coefs[9][108] = 16'h0000;
	mel_filter_coefs[9][109] = 16'h0000;
	mel_filter_coefs[9][110] = 16'h0000;
	mel_filter_coefs[9][111] = 16'h0000;
	mel_filter_coefs[9][112] = 16'h0000;
	mel_filter_coefs[9][113] = 16'h0000;
	mel_filter_coefs[9][114] = 16'h0000;
	mel_filter_coefs[9][115] = 16'h0000;
	mel_filter_coefs[9][116] = 16'h0000;
	mel_filter_coefs[9][117] = 16'h0000;
	mel_filter_coefs[9][118] = 16'h0000;
	mel_filter_coefs[9][119] = 16'h0000;
	mel_filter_coefs[9][120] = 16'h0000;
	mel_filter_coefs[9][121] = 16'h0000;
	mel_filter_coefs[9][122] = 16'h0000;
	mel_filter_coefs[9][123] = 16'h0000;
	mel_filter_coefs[9][124] = 16'h0000;
	mel_filter_coefs[9][125] = 16'h0000;
	mel_filter_coefs[9][126] = 16'h0000;
	mel_filter_coefs[9][127] = 16'h0000;
	mel_filter_coefs[9][128] = 16'h0000;
	mel_filter_coefs[9][129] = 16'h0000;
	mel_filter_coefs[9][130] = 16'h0000;
	mel_filter_coefs[9][131] = 16'h0000;
	mel_filter_coefs[9][132] = 16'h0000;
	mel_filter_coefs[9][133] = 16'h0000;
	mel_filter_coefs[9][134] = 16'h0000;
	mel_filter_coefs[9][135] = 16'h0000;
	mel_filter_coefs[9][136] = 16'h0000;
	mel_filter_coefs[9][137] = 16'h0000;
	mel_filter_coefs[9][138] = 16'h0000;
	mel_filter_coefs[9][139] = 16'h0000;
	mel_filter_coefs[9][140] = 16'h0000;
	mel_filter_coefs[9][141] = 16'h0000;
	mel_filter_coefs[9][142] = 16'h0000;
	mel_filter_coefs[9][143] = 16'h0000;
	mel_filter_coefs[9][144] = 16'h0000;
	mel_filter_coefs[9][145] = 16'h0000;
	mel_filter_coefs[9][146] = 16'h0000;
	mel_filter_coefs[9][147] = 16'h0000;
	mel_filter_coefs[9][148] = 16'h0000;
	mel_filter_coefs[9][149] = 16'h0000;
	mel_filter_coefs[9][150] = 16'h0000;
	mel_filter_coefs[9][151] = 16'h0000;
	mel_filter_coefs[9][152] = 16'h0000;
	mel_filter_coefs[9][153] = 16'h0000;
	mel_filter_coefs[9][154] = 16'h0000;
	mel_filter_coefs[9][155] = 16'h0000;
	mel_filter_coefs[9][156] = 16'h0000;
	mel_filter_coefs[9][157] = 16'h0000;
	mel_filter_coefs[9][158] = 16'h0000;
	mel_filter_coefs[9][159] = 16'h0000;
	mel_filter_coefs[9][160] = 16'h0000;
	mel_filter_coefs[9][161] = 16'h0000;
	mel_filter_coefs[9][162] = 16'h0000;
	mel_filter_coefs[9][163] = 16'h0000;
	mel_filter_coefs[9][164] = 16'h0000;
	mel_filter_coefs[9][165] = 16'h0000;
	mel_filter_coefs[9][166] = 16'h0000;
	mel_filter_coefs[9][167] = 16'h0000;
	mel_filter_coefs[9][168] = 16'h0000;
	mel_filter_coefs[9][169] = 16'h0000;
	mel_filter_coefs[9][170] = 16'h0000;
	mel_filter_coefs[9][171] = 16'h0000;
	mel_filter_coefs[9][172] = 16'h0000;
	mel_filter_coefs[9][173] = 16'h0000;
	mel_filter_coefs[9][174] = 16'h0000;
	mel_filter_coefs[9][175] = 16'h0000;
	mel_filter_coefs[9][176] = 16'h0000;
	mel_filter_coefs[9][177] = 16'h0000;
	mel_filter_coefs[9][178] = 16'h0000;
	mel_filter_coefs[9][179] = 16'h0000;
	mel_filter_coefs[9][180] = 16'h0000;
	mel_filter_coefs[9][181] = 16'h0000;
	mel_filter_coefs[9][182] = 16'h0000;
	mel_filter_coefs[9][183] = 16'h0000;
	mel_filter_coefs[9][184] = 16'h0000;
	mel_filter_coefs[9][185] = 16'h0000;
	mel_filter_coefs[9][186] = 16'h0000;
	mel_filter_coefs[9][187] = 16'h0000;
	mel_filter_coefs[9][188] = 16'h0000;
	mel_filter_coefs[9][189] = 16'h0000;
	mel_filter_coefs[9][190] = 16'h0000;
	mel_filter_coefs[9][191] = 16'h0000;
	mel_filter_coefs[9][192] = 16'h0000;
	mel_filter_coefs[9][193] = 16'h0000;
	mel_filter_coefs[9][194] = 16'h0000;
	mel_filter_coefs[9][195] = 16'h0000;
	mel_filter_coefs[9][196] = 16'h0000;
	mel_filter_coefs[9][197] = 16'h0000;
	mel_filter_coefs[9][198] = 16'h0000;
	mel_filter_coefs[9][199] = 16'h0000;
	mel_filter_coefs[9][200] = 16'h0000;
	mel_filter_coefs[9][201] = 16'h0000;
	mel_filter_coefs[9][202] = 16'h0000;
	mel_filter_coefs[9][203] = 16'h0000;
	mel_filter_coefs[9][204] = 16'h0000;
	mel_filter_coefs[9][205] = 16'h0000;
	mel_filter_coefs[9][206] = 16'h0000;
	mel_filter_coefs[9][207] = 16'h0000;
	mel_filter_coefs[9][208] = 16'h0000;
	mel_filter_coefs[9][209] = 16'h0000;
	mel_filter_coefs[9][210] = 16'h0000;
	mel_filter_coefs[9][211] = 16'h0000;
	mel_filter_coefs[9][212] = 16'h0000;
	mel_filter_coefs[9][213] = 16'h0000;
	mel_filter_coefs[9][214] = 16'h0000;
	mel_filter_coefs[9][215] = 16'h0000;
	mel_filter_coefs[9][216] = 16'h0000;
	mel_filter_coefs[9][217] = 16'h0000;
	mel_filter_coefs[9][218] = 16'h0000;
	mel_filter_coefs[9][219] = 16'h0000;
	mel_filter_coefs[9][220] = 16'h0000;
	mel_filter_coefs[9][221] = 16'h0000;
	mel_filter_coefs[9][222] = 16'h0000;
	mel_filter_coefs[9][223] = 16'h0000;
	mel_filter_coefs[9][224] = 16'h0000;
	mel_filter_coefs[9][225] = 16'h0000;
	mel_filter_coefs[9][226] = 16'h0000;
	mel_filter_coefs[9][227] = 16'h0000;
	mel_filter_coefs[9][228] = 16'h0000;
	mel_filter_coefs[9][229] = 16'h0000;
	mel_filter_coefs[9][230] = 16'h0000;
	mel_filter_coefs[9][231] = 16'h0000;
	mel_filter_coefs[9][232] = 16'h0000;
	mel_filter_coefs[9][233] = 16'h0000;
	mel_filter_coefs[9][234] = 16'h0000;
	mel_filter_coefs[9][235] = 16'h0000;
	mel_filter_coefs[9][236] = 16'h0000;
	mel_filter_coefs[9][237] = 16'h0000;
	mel_filter_coefs[9][238] = 16'h0000;
	mel_filter_coefs[9][239] = 16'h0000;
	mel_filter_coefs[9][240] = 16'h0000;
	mel_filter_coefs[9][241] = 16'h0000;
	mel_filter_coefs[9][242] = 16'h0000;
	mel_filter_coefs[9][243] = 16'h0000;
	mel_filter_coefs[9][244] = 16'h0000;
	mel_filter_coefs[9][245] = 16'h0000;
	mel_filter_coefs[9][246] = 16'h0000;
	mel_filter_coefs[9][247] = 16'h0000;
	mel_filter_coefs[9][248] = 16'h0000;
	mel_filter_coefs[9][249] = 16'h0000;
	mel_filter_coefs[9][250] = 16'h0000;
	mel_filter_coefs[9][251] = 16'h0000;
	mel_filter_coefs[9][252] = 16'h0000;
	mel_filter_coefs[9][253] = 16'h0000;
	mel_filter_coefs[9][254] = 16'h0000;
	mel_filter_coefs[9][255] = 16'h0000;
	mel_filter_coefs[10][0] = 16'h0000;
	mel_filter_coefs[10][1] = 16'h0000;
	mel_filter_coefs[10][2] = 16'h0000;
	mel_filter_coefs[10][3] = 16'h0000;
	mel_filter_coefs[10][4] = 16'h0000;
	mel_filter_coefs[10][5] = 16'h0000;
	mel_filter_coefs[10][6] = 16'h0000;
	mel_filter_coefs[10][7] = 16'h0000;
	mel_filter_coefs[10][8] = 16'h0000;
	mel_filter_coefs[10][9] = 16'h0000;
	mel_filter_coefs[10][10] = 16'h0000;
	mel_filter_coefs[10][11] = 16'h0000;
	mel_filter_coefs[10][12] = 16'h0000;
	mel_filter_coefs[10][13] = 16'h0000;
	mel_filter_coefs[10][14] = 16'h0000;
	mel_filter_coefs[10][15] = 16'h0000;
	mel_filter_coefs[10][16] = 16'h0000;
	mel_filter_coefs[10][17] = 16'h0000;
	mel_filter_coefs[10][18] = 16'h0000;
	mel_filter_coefs[10][19] = 16'h02CC;
	mel_filter_coefs[10][20] = 16'h33BE;
	mel_filter_coefs[10][21] = 16'h64AF;
	mel_filter_coefs[10][22] = 16'h6BA9;
	mel_filter_coefs[10][23] = 16'h3DA2;
	mel_filter_coefs[10][24] = 16'h0F9C;
	mel_filter_coefs[10][25] = 16'h0000;
	mel_filter_coefs[10][26] = 16'h0000;
	mel_filter_coefs[10][27] = 16'h0000;
	mel_filter_coefs[10][28] = 16'h0000;
	mel_filter_coefs[10][29] = 16'h0000;
	mel_filter_coefs[10][30] = 16'h0000;
	mel_filter_coefs[10][31] = 16'h0000;
	mel_filter_coefs[10][32] = 16'h0000;
	mel_filter_coefs[10][33] = 16'h0000;
	mel_filter_coefs[10][34] = 16'h0000;
	mel_filter_coefs[10][35] = 16'h0000;
	mel_filter_coefs[10][36] = 16'h0000;
	mel_filter_coefs[10][37] = 16'h0000;
	mel_filter_coefs[10][38] = 16'h0000;
	mel_filter_coefs[10][39] = 16'h0000;
	mel_filter_coefs[10][40] = 16'h0000;
	mel_filter_coefs[10][41] = 16'h0000;
	mel_filter_coefs[10][42] = 16'h0000;
	mel_filter_coefs[10][43] = 16'h0000;
	mel_filter_coefs[10][44] = 16'h0000;
	mel_filter_coefs[10][45] = 16'h0000;
	mel_filter_coefs[10][46] = 16'h0000;
	mel_filter_coefs[10][47] = 16'h0000;
	mel_filter_coefs[10][48] = 16'h0000;
	mel_filter_coefs[10][49] = 16'h0000;
	mel_filter_coefs[10][50] = 16'h0000;
	mel_filter_coefs[10][51] = 16'h0000;
	mel_filter_coefs[10][52] = 16'h0000;
	mel_filter_coefs[10][53] = 16'h0000;
	mel_filter_coefs[10][54] = 16'h0000;
	mel_filter_coefs[10][55] = 16'h0000;
	mel_filter_coefs[10][56] = 16'h0000;
	mel_filter_coefs[10][57] = 16'h0000;
	mel_filter_coefs[10][58] = 16'h0000;
	mel_filter_coefs[10][59] = 16'h0000;
	mel_filter_coefs[10][60] = 16'h0000;
	mel_filter_coefs[10][61] = 16'h0000;
	mel_filter_coefs[10][62] = 16'h0000;
	mel_filter_coefs[10][63] = 16'h0000;
	mel_filter_coefs[10][64] = 16'h0000;
	mel_filter_coefs[10][65] = 16'h0000;
	mel_filter_coefs[10][66] = 16'h0000;
	mel_filter_coefs[10][67] = 16'h0000;
	mel_filter_coefs[10][68] = 16'h0000;
	mel_filter_coefs[10][69] = 16'h0000;
	mel_filter_coefs[10][70] = 16'h0000;
	mel_filter_coefs[10][71] = 16'h0000;
	mel_filter_coefs[10][72] = 16'h0000;
	mel_filter_coefs[10][73] = 16'h0000;
	mel_filter_coefs[10][74] = 16'h0000;
	mel_filter_coefs[10][75] = 16'h0000;
	mel_filter_coefs[10][76] = 16'h0000;
	mel_filter_coefs[10][77] = 16'h0000;
	mel_filter_coefs[10][78] = 16'h0000;
	mel_filter_coefs[10][79] = 16'h0000;
	mel_filter_coefs[10][80] = 16'h0000;
	mel_filter_coefs[10][81] = 16'h0000;
	mel_filter_coefs[10][82] = 16'h0000;
	mel_filter_coefs[10][83] = 16'h0000;
	mel_filter_coefs[10][84] = 16'h0000;
	mel_filter_coefs[10][85] = 16'h0000;
	mel_filter_coefs[10][86] = 16'h0000;
	mel_filter_coefs[10][87] = 16'h0000;
	mel_filter_coefs[10][88] = 16'h0000;
	mel_filter_coefs[10][89] = 16'h0000;
	mel_filter_coefs[10][90] = 16'h0000;
	mel_filter_coefs[10][91] = 16'h0000;
	mel_filter_coefs[10][92] = 16'h0000;
	mel_filter_coefs[10][93] = 16'h0000;
	mel_filter_coefs[10][94] = 16'h0000;
	mel_filter_coefs[10][95] = 16'h0000;
	mel_filter_coefs[10][96] = 16'h0000;
	mel_filter_coefs[10][97] = 16'h0000;
	mel_filter_coefs[10][98] = 16'h0000;
	mel_filter_coefs[10][99] = 16'h0000;
	mel_filter_coefs[10][100] = 16'h0000;
	mel_filter_coefs[10][101] = 16'h0000;
	mel_filter_coefs[10][102] = 16'h0000;
	mel_filter_coefs[10][103] = 16'h0000;
	mel_filter_coefs[10][104] = 16'h0000;
	mel_filter_coefs[10][105] = 16'h0000;
	mel_filter_coefs[10][106] = 16'h0000;
	mel_filter_coefs[10][107] = 16'h0000;
	mel_filter_coefs[10][108] = 16'h0000;
	mel_filter_coefs[10][109] = 16'h0000;
	mel_filter_coefs[10][110] = 16'h0000;
	mel_filter_coefs[10][111] = 16'h0000;
	mel_filter_coefs[10][112] = 16'h0000;
	mel_filter_coefs[10][113] = 16'h0000;
	mel_filter_coefs[10][114] = 16'h0000;
	mel_filter_coefs[10][115] = 16'h0000;
	mel_filter_coefs[10][116] = 16'h0000;
	mel_filter_coefs[10][117] = 16'h0000;
	mel_filter_coefs[10][118] = 16'h0000;
	mel_filter_coefs[10][119] = 16'h0000;
	mel_filter_coefs[10][120] = 16'h0000;
	mel_filter_coefs[10][121] = 16'h0000;
	mel_filter_coefs[10][122] = 16'h0000;
	mel_filter_coefs[10][123] = 16'h0000;
	mel_filter_coefs[10][124] = 16'h0000;
	mel_filter_coefs[10][125] = 16'h0000;
	mel_filter_coefs[10][126] = 16'h0000;
	mel_filter_coefs[10][127] = 16'h0000;
	mel_filter_coefs[10][128] = 16'h0000;
	mel_filter_coefs[10][129] = 16'h0000;
	mel_filter_coefs[10][130] = 16'h0000;
	mel_filter_coefs[10][131] = 16'h0000;
	mel_filter_coefs[10][132] = 16'h0000;
	mel_filter_coefs[10][133] = 16'h0000;
	mel_filter_coefs[10][134] = 16'h0000;
	mel_filter_coefs[10][135] = 16'h0000;
	mel_filter_coefs[10][136] = 16'h0000;
	mel_filter_coefs[10][137] = 16'h0000;
	mel_filter_coefs[10][138] = 16'h0000;
	mel_filter_coefs[10][139] = 16'h0000;
	mel_filter_coefs[10][140] = 16'h0000;
	mel_filter_coefs[10][141] = 16'h0000;
	mel_filter_coefs[10][142] = 16'h0000;
	mel_filter_coefs[10][143] = 16'h0000;
	mel_filter_coefs[10][144] = 16'h0000;
	mel_filter_coefs[10][145] = 16'h0000;
	mel_filter_coefs[10][146] = 16'h0000;
	mel_filter_coefs[10][147] = 16'h0000;
	mel_filter_coefs[10][148] = 16'h0000;
	mel_filter_coefs[10][149] = 16'h0000;
	mel_filter_coefs[10][150] = 16'h0000;
	mel_filter_coefs[10][151] = 16'h0000;
	mel_filter_coefs[10][152] = 16'h0000;
	mel_filter_coefs[10][153] = 16'h0000;
	mel_filter_coefs[10][154] = 16'h0000;
	mel_filter_coefs[10][155] = 16'h0000;
	mel_filter_coefs[10][156] = 16'h0000;
	mel_filter_coefs[10][157] = 16'h0000;
	mel_filter_coefs[10][158] = 16'h0000;
	mel_filter_coefs[10][159] = 16'h0000;
	mel_filter_coefs[10][160] = 16'h0000;
	mel_filter_coefs[10][161] = 16'h0000;
	mel_filter_coefs[10][162] = 16'h0000;
	mel_filter_coefs[10][163] = 16'h0000;
	mel_filter_coefs[10][164] = 16'h0000;
	mel_filter_coefs[10][165] = 16'h0000;
	mel_filter_coefs[10][166] = 16'h0000;
	mel_filter_coefs[10][167] = 16'h0000;
	mel_filter_coefs[10][168] = 16'h0000;
	mel_filter_coefs[10][169] = 16'h0000;
	mel_filter_coefs[10][170] = 16'h0000;
	mel_filter_coefs[10][171] = 16'h0000;
	mel_filter_coefs[10][172] = 16'h0000;
	mel_filter_coefs[10][173] = 16'h0000;
	mel_filter_coefs[10][174] = 16'h0000;
	mel_filter_coefs[10][175] = 16'h0000;
	mel_filter_coefs[10][176] = 16'h0000;
	mel_filter_coefs[10][177] = 16'h0000;
	mel_filter_coefs[10][178] = 16'h0000;
	mel_filter_coefs[10][179] = 16'h0000;
	mel_filter_coefs[10][180] = 16'h0000;
	mel_filter_coefs[10][181] = 16'h0000;
	mel_filter_coefs[10][182] = 16'h0000;
	mel_filter_coefs[10][183] = 16'h0000;
	mel_filter_coefs[10][184] = 16'h0000;
	mel_filter_coefs[10][185] = 16'h0000;
	mel_filter_coefs[10][186] = 16'h0000;
	mel_filter_coefs[10][187] = 16'h0000;
	mel_filter_coefs[10][188] = 16'h0000;
	mel_filter_coefs[10][189] = 16'h0000;
	mel_filter_coefs[10][190] = 16'h0000;
	mel_filter_coefs[10][191] = 16'h0000;
	mel_filter_coefs[10][192] = 16'h0000;
	mel_filter_coefs[10][193] = 16'h0000;
	mel_filter_coefs[10][194] = 16'h0000;
	mel_filter_coefs[10][195] = 16'h0000;
	mel_filter_coefs[10][196] = 16'h0000;
	mel_filter_coefs[10][197] = 16'h0000;
	mel_filter_coefs[10][198] = 16'h0000;
	mel_filter_coefs[10][199] = 16'h0000;
	mel_filter_coefs[10][200] = 16'h0000;
	mel_filter_coefs[10][201] = 16'h0000;
	mel_filter_coefs[10][202] = 16'h0000;
	mel_filter_coefs[10][203] = 16'h0000;
	mel_filter_coefs[10][204] = 16'h0000;
	mel_filter_coefs[10][205] = 16'h0000;
	mel_filter_coefs[10][206] = 16'h0000;
	mel_filter_coefs[10][207] = 16'h0000;
	mel_filter_coefs[10][208] = 16'h0000;
	mel_filter_coefs[10][209] = 16'h0000;
	mel_filter_coefs[10][210] = 16'h0000;
	mel_filter_coefs[10][211] = 16'h0000;
	mel_filter_coefs[10][212] = 16'h0000;
	mel_filter_coefs[10][213] = 16'h0000;
	mel_filter_coefs[10][214] = 16'h0000;
	mel_filter_coefs[10][215] = 16'h0000;
	mel_filter_coefs[10][216] = 16'h0000;
	mel_filter_coefs[10][217] = 16'h0000;
	mel_filter_coefs[10][218] = 16'h0000;
	mel_filter_coefs[10][219] = 16'h0000;
	mel_filter_coefs[10][220] = 16'h0000;
	mel_filter_coefs[10][221] = 16'h0000;
	mel_filter_coefs[10][222] = 16'h0000;
	mel_filter_coefs[10][223] = 16'h0000;
	mel_filter_coefs[10][224] = 16'h0000;
	mel_filter_coefs[10][225] = 16'h0000;
	mel_filter_coefs[10][226] = 16'h0000;
	mel_filter_coefs[10][227] = 16'h0000;
	mel_filter_coefs[10][228] = 16'h0000;
	mel_filter_coefs[10][229] = 16'h0000;
	mel_filter_coefs[10][230] = 16'h0000;
	mel_filter_coefs[10][231] = 16'h0000;
	mel_filter_coefs[10][232] = 16'h0000;
	mel_filter_coefs[10][233] = 16'h0000;
	mel_filter_coefs[10][234] = 16'h0000;
	mel_filter_coefs[10][235] = 16'h0000;
	mel_filter_coefs[10][236] = 16'h0000;
	mel_filter_coefs[10][237] = 16'h0000;
	mel_filter_coefs[10][238] = 16'h0000;
	mel_filter_coefs[10][239] = 16'h0000;
	mel_filter_coefs[10][240] = 16'h0000;
	mel_filter_coefs[10][241] = 16'h0000;
	mel_filter_coefs[10][242] = 16'h0000;
	mel_filter_coefs[10][243] = 16'h0000;
	mel_filter_coefs[10][244] = 16'h0000;
	mel_filter_coefs[10][245] = 16'h0000;
	mel_filter_coefs[10][246] = 16'h0000;
	mel_filter_coefs[10][247] = 16'h0000;
	mel_filter_coefs[10][248] = 16'h0000;
	mel_filter_coefs[10][249] = 16'h0000;
	mel_filter_coefs[10][250] = 16'h0000;
	mel_filter_coefs[10][251] = 16'h0000;
	mel_filter_coefs[10][252] = 16'h0000;
	mel_filter_coefs[10][253] = 16'h0000;
	mel_filter_coefs[10][254] = 16'h0000;
	mel_filter_coefs[10][255] = 16'h0000;
	mel_filter_coefs[11][0] = 16'h0000;
	mel_filter_coefs[11][1] = 16'h0000;
	mel_filter_coefs[11][2] = 16'h0000;
	mel_filter_coefs[11][3] = 16'h0000;
	mel_filter_coefs[11][4] = 16'h0000;
	mel_filter_coefs[11][5] = 16'h0000;
	mel_filter_coefs[11][6] = 16'h0000;
	mel_filter_coefs[11][7] = 16'h0000;
	mel_filter_coefs[11][8] = 16'h0000;
	mel_filter_coefs[11][9] = 16'h0000;
	mel_filter_coefs[11][10] = 16'h0000;
	mel_filter_coefs[11][11] = 16'h0000;
	mel_filter_coefs[11][12] = 16'h0000;
	mel_filter_coefs[11][13] = 16'h0000;
	mel_filter_coefs[11][14] = 16'h0000;
	mel_filter_coefs[11][15] = 16'h0000;
	mel_filter_coefs[11][16] = 16'h0000;
	mel_filter_coefs[11][17] = 16'h0000;
	mel_filter_coefs[11][18] = 16'h0000;
	mel_filter_coefs[11][19] = 16'h0000;
	mel_filter_coefs[11][20] = 16'h0000;
	mel_filter_coefs[11][21] = 16'h0000;
	mel_filter_coefs[11][22] = 16'h1457;
	mel_filter_coefs[11][23] = 16'h425E;
	mel_filter_coefs[11][24] = 16'h7064;
	mel_filter_coefs[11][25] = 16'h6365;
	mel_filter_coefs[11][26] = 16'h381D;
	mel_filter_coefs[11][27] = 16'h0CD5;
	mel_filter_coefs[11][28] = 16'h0000;
	mel_filter_coefs[11][29] = 16'h0000;
	mel_filter_coefs[11][30] = 16'h0000;
	mel_filter_coefs[11][31] = 16'h0000;
	mel_filter_coefs[11][32] = 16'h0000;
	mel_filter_coefs[11][33] = 16'h0000;
	mel_filter_coefs[11][34] = 16'h0000;
	mel_filter_coefs[11][35] = 16'h0000;
	mel_filter_coefs[11][36] = 16'h0000;
	mel_filter_coefs[11][37] = 16'h0000;
	mel_filter_coefs[11][38] = 16'h0000;
	mel_filter_coefs[11][39] = 16'h0000;
	mel_filter_coefs[11][40] = 16'h0000;
	mel_filter_coefs[11][41] = 16'h0000;
	mel_filter_coefs[11][42] = 16'h0000;
	mel_filter_coefs[11][43] = 16'h0000;
	mel_filter_coefs[11][44] = 16'h0000;
	mel_filter_coefs[11][45] = 16'h0000;
	mel_filter_coefs[11][46] = 16'h0000;
	mel_filter_coefs[11][47] = 16'h0000;
	mel_filter_coefs[11][48] = 16'h0000;
	mel_filter_coefs[11][49] = 16'h0000;
	mel_filter_coefs[11][50] = 16'h0000;
	mel_filter_coefs[11][51] = 16'h0000;
	mel_filter_coefs[11][52] = 16'h0000;
	mel_filter_coefs[11][53] = 16'h0000;
	mel_filter_coefs[11][54] = 16'h0000;
	mel_filter_coefs[11][55] = 16'h0000;
	mel_filter_coefs[11][56] = 16'h0000;
	mel_filter_coefs[11][57] = 16'h0000;
	mel_filter_coefs[11][58] = 16'h0000;
	mel_filter_coefs[11][59] = 16'h0000;
	mel_filter_coefs[11][60] = 16'h0000;
	mel_filter_coefs[11][61] = 16'h0000;
	mel_filter_coefs[11][62] = 16'h0000;
	mel_filter_coefs[11][63] = 16'h0000;
	mel_filter_coefs[11][64] = 16'h0000;
	mel_filter_coefs[11][65] = 16'h0000;
	mel_filter_coefs[11][66] = 16'h0000;
	mel_filter_coefs[11][67] = 16'h0000;
	mel_filter_coefs[11][68] = 16'h0000;
	mel_filter_coefs[11][69] = 16'h0000;
	mel_filter_coefs[11][70] = 16'h0000;
	mel_filter_coefs[11][71] = 16'h0000;
	mel_filter_coefs[11][72] = 16'h0000;
	mel_filter_coefs[11][73] = 16'h0000;
	mel_filter_coefs[11][74] = 16'h0000;
	mel_filter_coefs[11][75] = 16'h0000;
	mel_filter_coefs[11][76] = 16'h0000;
	mel_filter_coefs[11][77] = 16'h0000;
	mel_filter_coefs[11][78] = 16'h0000;
	mel_filter_coefs[11][79] = 16'h0000;
	mel_filter_coefs[11][80] = 16'h0000;
	mel_filter_coefs[11][81] = 16'h0000;
	mel_filter_coefs[11][82] = 16'h0000;
	mel_filter_coefs[11][83] = 16'h0000;
	mel_filter_coefs[11][84] = 16'h0000;
	mel_filter_coefs[11][85] = 16'h0000;
	mel_filter_coefs[11][86] = 16'h0000;
	mel_filter_coefs[11][87] = 16'h0000;
	mel_filter_coefs[11][88] = 16'h0000;
	mel_filter_coefs[11][89] = 16'h0000;
	mel_filter_coefs[11][90] = 16'h0000;
	mel_filter_coefs[11][91] = 16'h0000;
	mel_filter_coefs[11][92] = 16'h0000;
	mel_filter_coefs[11][93] = 16'h0000;
	mel_filter_coefs[11][94] = 16'h0000;
	mel_filter_coefs[11][95] = 16'h0000;
	mel_filter_coefs[11][96] = 16'h0000;
	mel_filter_coefs[11][97] = 16'h0000;
	mel_filter_coefs[11][98] = 16'h0000;
	mel_filter_coefs[11][99] = 16'h0000;
	mel_filter_coefs[11][100] = 16'h0000;
	mel_filter_coefs[11][101] = 16'h0000;
	mel_filter_coefs[11][102] = 16'h0000;
	mel_filter_coefs[11][103] = 16'h0000;
	mel_filter_coefs[11][104] = 16'h0000;
	mel_filter_coefs[11][105] = 16'h0000;
	mel_filter_coefs[11][106] = 16'h0000;
	mel_filter_coefs[11][107] = 16'h0000;
	mel_filter_coefs[11][108] = 16'h0000;
	mel_filter_coefs[11][109] = 16'h0000;
	mel_filter_coefs[11][110] = 16'h0000;
	mel_filter_coefs[11][111] = 16'h0000;
	mel_filter_coefs[11][112] = 16'h0000;
	mel_filter_coefs[11][113] = 16'h0000;
	mel_filter_coefs[11][114] = 16'h0000;
	mel_filter_coefs[11][115] = 16'h0000;
	mel_filter_coefs[11][116] = 16'h0000;
	mel_filter_coefs[11][117] = 16'h0000;
	mel_filter_coefs[11][118] = 16'h0000;
	mel_filter_coefs[11][119] = 16'h0000;
	mel_filter_coefs[11][120] = 16'h0000;
	mel_filter_coefs[11][121] = 16'h0000;
	mel_filter_coefs[11][122] = 16'h0000;
	mel_filter_coefs[11][123] = 16'h0000;
	mel_filter_coefs[11][124] = 16'h0000;
	mel_filter_coefs[11][125] = 16'h0000;
	mel_filter_coefs[11][126] = 16'h0000;
	mel_filter_coefs[11][127] = 16'h0000;
	mel_filter_coefs[11][128] = 16'h0000;
	mel_filter_coefs[11][129] = 16'h0000;
	mel_filter_coefs[11][130] = 16'h0000;
	mel_filter_coefs[11][131] = 16'h0000;
	mel_filter_coefs[11][132] = 16'h0000;
	mel_filter_coefs[11][133] = 16'h0000;
	mel_filter_coefs[11][134] = 16'h0000;
	mel_filter_coefs[11][135] = 16'h0000;
	mel_filter_coefs[11][136] = 16'h0000;
	mel_filter_coefs[11][137] = 16'h0000;
	mel_filter_coefs[11][138] = 16'h0000;
	mel_filter_coefs[11][139] = 16'h0000;
	mel_filter_coefs[11][140] = 16'h0000;
	mel_filter_coefs[11][141] = 16'h0000;
	mel_filter_coefs[11][142] = 16'h0000;
	mel_filter_coefs[11][143] = 16'h0000;
	mel_filter_coefs[11][144] = 16'h0000;
	mel_filter_coefs[11][145] = 16'h0000;
	mel_filter_coefs[11][146] = 16'h0000;
	mel_filter_coefs[11][147] = 16'h0000;
	mel_filter_coefs[11][148] = 16'h0000;
	mel_filter_coefs[11][149] = 16'h0000;
	mel_filter_coefs[11][150] = 16'h0000;
	mel_filter_coefs[11][151] = 16'h0000;
	mel_filter_coefs[11][152] = 16'h0000;
	mel_filter_coefs[11][153] = 16'h0000;
	mel_filter_coefs[11][154] = 16'h0000;
	mel_filter_coefs[11][155] = 16'h0000;
	mel_filter_coefs[11][156] = 16'h0000;
	mel_filter_coefs[11][157] = 16'h0000;
	mel_filter_coefs[11][158] = 16'h0000;
	mel_filter_coefs[11][159] = 16'h0000;
	mel_filter_coefs[11][160] = 16'h0000;
	mel_filter_coefs[11][161] = 16'h0000;
	mel_filter_coefs[11][162] = 16'h0000;
	mel_filter_coefs[11][163] = 16'h0000;
	mel_filter_coefs[11][164] = 16'h0000;
	mel_filter_coefs[11][165] = 16'h0000;
	mel_filter_coefs[11][166] = 16'h0000;
	mel_filter_coefs[11][167] = 16'h0000;
	mel_filter_coefs[11][168] = 16'h0000;
	mel_filter_coefs[11][169] = 16'h0000;
	mel_filter_coefs[11][170] = 16'h0000;
	mel_filter_coefs[11][171] = 16'h0000;
	mel_filter_coefs[11][172] = 16'h0000;
	mel_filter_coefs[11][173] = 16'h0000;
	mel_filter_coefs[11][174] = 16'h0000;
	mel_filter_coefs[11][175] = 16'h0000;
	mel_filter_coefs[11][176] = 16'h0000;
	mel_filter_coefs[11][177] = 16'h0000;
	mel_filter_coefs[11][178] = 16'h0000;
	mel_filter_coefs[11][179] = 16'h0000;
	mel_filter_coefs[11][180] = 16'h0000;
	mel_filter_coefs[11][181] = 16'h0000;
	mel_filter_coefs[11][182] = 16'h0000;
	mel_filter_coefs[11][183] = 16'h0000;
	mel_filter_coefs[11][184] = 16'h0000;
	mel_filter_coefs[11][185] = 16'h0000;
	mel_filter_coefs[11][186] = 16'h0000;
	mel_filter_coefs[11][187] = 16'h0000;
	mel_filter_coefs[11][188] = 16'h0000;
	mel_filter_coefs[11][189] = 16'h0000;
	mel_filter_coefs[11][190] = 16'h0000;
	mel_filter_coefs[11][191] = 16'h0000;
	mel_filter_coefs[11][192] = 16'h0000;
	mel_filter_coefs[11][193] = 16'h0000;
	mel_filter_coefs[11][194] = 16'h0000;
	mel_filter_coefs[11][195] = 16'h0000;
	mel_filter_coefs[11][196] = 16'h0000;
	mel_filter_coefs[11][197] = 16'h0000;
	mel_filter_coefs[11][198] = 16'h0000;
	mel_filter_coefs[11][199] = 16'h0000;
	mel_filter_coefs[11][200] = 16'h0000;
	mel_filter_coefs[11][201] = 16'h0000;
	mel_filter_coefs[11][202] = 16'h0000;
	mel_filter_coefs[11][203] = 16'h0000;
	mel_filter_coefs[11][204] = 16'h0000;
	mel_filter_coefs[11][205] = 16'h0000;
	mel_filter_coefs[11][206] = 16'h0000;
	mel_filter_coefs[11][207] = 16'h0000;
	mel_filter_coefs[11][208] = 16'h0000;
	mel_filter_coefs[11][209] = 16'h0000;
	mel_filter_coefs[11][210] = 16'h0000;
	mel_filter_coefs[11][211] = 16'h0000;
	mel_filter_coefs[11][212] = 16'h0000;
	mel_filter_coefs[11][213] = 16'h0000;
	mel_filter_coefs[11][214] = 16'h0000;
	mel_filter_coefs[11][215] = 16'h0000;
	mel_filter_coefs[11][216] = 16'h0000;
	mel_filter_coefs[11][217] = 16'h0000;
	mel_filter_coefs[11][218] = 16'h0000;
	mel_filter_coefs[11][219] = 16'h0000;
	mel_filter_coefs[11][220] = 16'h0000;
	mel_filter_coefs[11][221] = 16'h0000;
	mel_filter_coefs[11][222] = 16'h0000;
	mel_filter_coefs[11][223] = 16'h0000;
	mel_filter_coefs[11][224] = 16'h0000;
	mel_filter_coefs[11][225] = 16'h0000;
	mel_filter_coefs[11][226] = 16'h0000;
	mel_filter_coefs[11][227] = 16'h0000;
	mel_filter_coefs[11][228] = 16'h0000;
	mel_filter_coefs[11][229] = 16'h0000;
	mel_filter_coefs[11][230] = 16'h0000;
	mel_filter_coefs[11][231] = 16'h0000;
	mel_filter_coefs[11][232] = 16'h0000;
	mel_filter_coefs[11][233] = 16'h0000;
	mel_filter_coefs[11][234] = 16'h0000;
	mel_filter_coefs[11][235] = 16'h0000;
	mel_filter_coefs[11][236] = 16'h0000;
	mel_filter_coefs[11][237] = 16'h0000;
	mel_filter_coefs[11][238] = 16'h0000;
	mel_filter_coefs[11][239] = 16'h0000;
	mel_filter_coefs[11][240] = 16'h0000;
	mel_filter_coefs[11][241] = 16'h0000;
	mel_filter_coefs[11][242] = 16'h0000;
	mel_filter_coefs[11][243] = 16'h0000;
	mel_filter_coefs[11][244] = 16'h0000;
	mel_filter_coefs[11][245] = 16'h0000;
	mel_filter_coefs[11][246] = 16'h0000;
	mel_filter_coefs[11][247] = 16'h0000;
	mel_filter_coefs[11][248] = 16'h0000;
	mel_filter_coefs[11][249] = 16'h0000;
	mel_filter_coefs[11][250] = 16'h0000;
	mel_filter_coefs[11][251] = 16'h0000;
	mel_filter_coefs[11][252] = 16'h0000;
	mel_filter_coefs[11][253] = 16'h0000;
	mel_filter_coefs[11][254] = 16'h0000;
	mel_filter_coefs[11][255] = 16'h0000;
	mel_filter_coefs[12][0] = 16'h0000;
	mel_filter_coefs[12][1] = 16'h0000;
	mel_filter_coefs[12][2] = 16'h0000;
	mel_filter_coefs[12][3] = 16'h0000;
	mel_filter_coefs[12][4] = 16'h0000;
	mel_filter_coefs[12][5] = 16'h0000;
	mel_filter_coefs[12][6] = 16'h0000;
	mel_filter_coefs[12][7] = 16'h0000;
	mel_filter_coefs[12][8] = 16'h0000;
	mel_filter_coefs[12][9] = 16'h0000;
	mel_filter_coefs[12][10] = 16'h0000;
	mel_filter_coefs[12][11] = 16'h0000;
	mel_filter_coefs[12][12] = 16'h0000;
	mel_filter_coefs[12][13] = 16'h0000;
	mel_filter_coefs[12][14] = 16'h0000;
	mel_filter_coefs[12][15] = 16'h0000;
	mel_filter_coefs[12][16] = 16'h0000;
	mel_filter_coefs[12][17] = 16'h0000;
	mel_filter_coefs[12][18] = 16'h0000;
	mel_filter_coefs[12][19] = 16'h0000;
	mel_filter_coefs[12][20] = 16'h0000;
	mel_filter_coefs[12][21] = 16'h0000;
	mel_filter_coefs[12][22] = 16'h0000;
	mel_filter_coefs[12][23] = 16'h0000;
	mel_filter_coefs[12][24] = 16'h0000;
	mel_filter_coefs[12][25] = 16'h1C9B;
	mel_filter_coefs[12][26] = 16'h47E3;
	mel_filter_coefs[12][27] = 16'h732B;
	mel_filter_coefs[12][28] = 16'h635D;
	mel_filter_coefs[12][29] = 16'h3AA9;
	mel_filter_coefs[12][30] = 16'h11F5;
	mel_filter_coefs[12][31] = 16'h0000;
	mel_filter_coefs[12][32] = 16'h0000;
	mel_filter_coefs[12][33] = 16'h0000;
	mel_filter_coefs[12][34] = 16'h0000;
	mel_filter_coefs[12][35] = 16'h0000;
	mel_filter_coefs[12][36] = 16'h0000;
	mel_filter_coefs[12][37] = 16'h0000;
	mel_filter_coefs[12][38] = 16'h0000;
	mel_filter_coefs[12][39] = 16'h0000;
	mel_filter_coefs[12][40] = 16'h0000;
	mel_filter_coefs[12][41] = 16'h0000;
	mel_filter_coefs[12][42] = 16'h0000;
	mel_filter_coefs[12][43] = 16'h0000;
	mel_filter_coefs[12][44] = 16'h0000;
	mel_filter_coefs[12][45] = 16'h0000;
	mel_filter_coefs[12][46] = 16'h0000;
	mel_filter_coefs[12][47] = 16'h0000;
	mel_filter_coefs[12][48] = 16'h0000;
	mel_filter_coefs[12][49] = 16'h0000;
	mel_filter_coefs[12][50] = 16'h0000;
	mel_filter_coefs[12][51] = 16'h0000;
	mel_filter_coefs[12][52] = 16'h0000;
	mel_filter_coefs[12][53] = 16'h0000;
	mel_filter_coefs[12][54] = 16'h0000;
	mel_filter_coefs[12][55] = 16'h0000;
	mel_filter_coefs[12][56] = 16'h0000;
	mel_filter_coefs[12][57] = 16'h0000;
	mel_filter_coefs[12][58] = 16'h0000;
	mel_filter_coefs[12][59] = 16'h0000;
	mel_filter_coefs[12][60] = 16'h0000;
	mel_filter_coefs[12][61] = 16'h0000;
	mel_filter_coefs[12][62] = 16'h0000;
	mel_filter_coefs[12][63] = 16'h0000;
	mel_filter_coefs[12][64] = 16'h0000;
	mel_filter_coefs[12][65] = 16'h0000;
	mel_filter_coefs[12][66] = 16'h0000;
	mel_filter_coefs[12][67] = 16'h0000;
	mel_filter_coefs[12][68] = 16'h0000;
	mel_filter_coefs[12][69] = 16'h0000;
	mel_filter_coefs[12][70] = 16'h0000;
	mel_filter_coefs[12][71] = 16'h0000;
	mel_filter_coefs[12][72] = 16'h0000;
	mel_filter_coefs[12][73] = 16'h0000;
	mel_filter_coefs[12][74] = 16'h0000;
	mel_filter_coefs[12][75] = 16'h0000;
	mel_filter_coefs[12][76] = 16'h0000;
	mel_filter_coefs[12][77] = 16'h0000;
	mel_filter_coefs[12][78] = 16'h0000;
	mel_filter_coefs[12][79] = 16'h0000;
	mel_filter_coefs[12][80] = 16'h0000;
	mel_filter_coefs[12][81] = 16'h0000;
	mel_filter_coefs[12][82] = 16'h0000;
	mel_filter_coefs[12][83] = 16'h0000;
	mel_filter_coefs[12][84] = 16'h0000;
	mel_filter_coefs[12][85] = 16'h0000;
	mel_filter_coefs[12][86] = 16'h0000;
	mel_filter_coefs[12][87] = 16'h0000;
	mel_filter_coefs[12][88] = 16'h0000;
	mel_filter_coefs[12][89] = 16'h0000;
	mel_filter_coefs[12][90] = 16'h0000;
	mel_filter_coefs[12][91] = 16'h0000;
	mel_filter_coefs[12][92] = 16'h0000;
	mel_filter_coefs[12][93] = 16'h0000;
	mel_filter_coefs[12][94] = 16'h0000;
	mel_filter_coefs[12][95] = 16'h0000;
	mel_filter_coefs[12][96] = 16'h0000;
	mel_filter_coefs[12][97] = 16'h0000;
	mel_filter_coefs[12][98] = 16'h0000;
	mel_filter_coefs[12][99] = 16'h0000;
	mel_filter_coefs[12][100] = 16'h0000;
	mel_filter_coefs[12][101] = 16'h0000;
	mel_filter_coefs[12][102] = 16'h0000;
	mel_filter_coefs[12][103] = 16'h0000;
	mel_filter_coefs[12][104] = 16'h0000;
	mel_filter_coefs[12][105] = 16'h0000;
	mel_filter_coefs[12][106] = 16'h0000;
	mel_filter_coefs[12][107] = 16'h0000;
	mel_filter_coefs[12][108] = 16'h0000;
	mel_filter_coefs[12][109] = 16'h0000;
	mel_filter_coefs[12][110] = 16'h0000;
	mel_filter_coefs[12][111] = 16'h0000;
	mel_filter_coefs[12][112] = 16'h0000;
	mel_filter_coefs[12][113] = 16'h0000;
	mel_filter_coefs[12][114] = 16'h0000;
	mel_filter_coefs[12][115] = 16'h0000;
	mel_filter_coefs[12][116] = 16'h0000;
	mel_filter_coefs[12][117] = 16'h0000;
	mel_filter_coefs[12][118] = 16'h0000;
	mel_filter_coefs[12][119] = 16'h0000;
	mel_filter_coefs[12][120] = 16'h0000;
	mel_filter_coefs[12][121] = 16'h0000;
	mel_filter_coefs[12][122] = 16'h0000;
	mel_filter_coefs[12][123] = 16'h0000;
	mel_filter_coefs[12][124] = 16'h0000;
	mel_filter_coefs[12][125] = 16'h0000;
	mel_filter_coefs[12][126] = 16'h0000;
	mel_filter_coefs[12][127] = 16'h0000;
	mel_filter_coefs[12][128] = 16'h0000;
	mel_filter_coefs[12][129] = 16'h0000;
	mel_filter_coefs[12][130] = 16'h0000;
	mel_filter_coefs[12][131] = 16'h0000;
	mel_filter_coefs[12][132] = 16'h0000;
	mel_filter_coefs[12][133] = 16'h0000;
	mel_filter_coefs[12][134] = 16'h0000;
	mel_filter_coefs[12][135] = 16'h0000;
	mel_filter_coefs[12][136] = 16'h0000;
	mel_filter_coefs[12][137] = 16'h0000;
	mel_filter_coefs[12][138] = 16'h0000;
	mel_filter_coefs[12][139] = 16'h0000;
	mel_filter_coefs[12][140] = 16'h0000;
	mel_filter_coefs[12][141] = 16'h0000;
	mel_filter_coefs[12][142] = 16'h0000;
	mel_filter_coefs[12][143] = 16'h0000;
	mel_filter_coefs[12][144] = 16'h0000;
	mel_filter_coefs[12][145] = 16'h0000;
	mel_filter_coefs[12][146] = 16'h0000;
	mel_filter_coefs[12][147] = 16'h0000;
	mel_filter_coefs[12][148] = 16'h0000;
	mel_filter_coefs[12][149] = 16'h0000;
	mel_filter_coefs[12][150] = 16'h0000;
	mel_filter_coefs[12][151] = 16'h0000;
	mel_filter_coefs[12][152] = 16'h0000;
	mel_filter_coefs[12][153] = 16'h0000;
	mel_filter_coefs[12][154] = 16'h0000;
	mel_filter_coefs[12][155] = 16'h0000;
	mel_filter_coefs[12][156] = 16'h0000;
	mel_filter_coefs[12][157] = 16'h0000;
	mel_filter_coefs[12][158] = 16'h0000;
	mel_filter_coefs[12][159] = 16'h0000;
	mel_filter_coefs[12][160] = 16'h0000;
	mel_filter_coefs[12][161] = 16'h0000;
	mel_filter_coefs[12][162] = 16'h0000;
	mel_filter_coefs[12][163] = 16'h0000;
	mel_filter_coefs[12][164] = 16'h0000;
	mel_filter_coefs[12][165] = 16'h0000;
	mel_filter_coefs[12][166] = 16'h0000;
	mel_filter_coefs[12][167] = 16'h0000;
	mel_filter_coefs[12][168] = 16'h0000;
	mel_filter_coefs[12][169] = 16'h0000;
	mel_filter_coefs[12][170] = 16'h0000;
	mel_filter_coefs[12][171] = 16'h0000;
	mel_filter_coefs[12][172] = 16'h0000;
	mel_filter_coefs[12][173] = 16'h0000;
	mel_filter_coefs[12][174] = 16'h0000;
	mel_filter_coefs[12][175] = 16'h0000;
	mel_filter_coefs[12][176] = 16'h0000;
	mel_filter_coefs[12][177] = 16'h0000;
	mel_filter_coefs[12][178] = 16'h0000;
	mel_filter_coefs[12][179] = 16'h0000;
	mel_filter_coefs[12][180] = 16'h0000;
	mel_filter_coefs[12][181] = 16'h0000;
	mel_filter_coefs[12][182] = 16'h0000;
	mel_filter_coefs[12][183] = 16'h0000;
	mel_filter_coefs[12][184] = 16'h0000;
	mel_filter_coefs[12][185] = 16'h0000;
	mel_filter_coefs[12][186] = 16'h0000;
	mel_filter_coefs[12][187] = 16'h0000;
	mel_filter_coefs[12][188] = 16'h0000;
	mel_filter_coefs[12][189] = 16'h0000;
	mel_filter_coefs[12][190] = 16'h0000;
	mel_filter_coefs[12][191] = 16'h0000;
	mel_filter_coefs[12][192] = 16'h0000;
	mel_filter_coefs[12][193] = 16'h0000;
	mel_filter_coefs[12][194] = 16'h0000;
	mel_filter_coefs[12][195] = 16'h0000;
	mel_filter_coefs[12][196] = 16'h0000;
	mel_filter_coefs[12][197] = 16'h0000;
	mel_filter_coefs[12][198] = 16'h0000;
	mel_filter_coefs[12][199] = 16'h0000;
	mel_filter_coefs[12][200] = 16'h0000;
	mel_filter_coefs[12][201] = 16'h0000;
	mel_filter_coefs[12][202] = 16'h0000;
	mel_filter_coefs[12][203] = 16'h0000;
	mel_filter_coefs[12][204] = 16'h0000;
	mel_filter_coefs[12][205] = 16'h0000;
	mel_filter_coefs[12][206] = 16'h0000;
	mel_filter_coefs[12][207] = 16'h0000;
	mel_filter_coefs[12][208] = 16'h0000;
	mel_filter_coefs[12][209] = 16'h0000;
	mel_filter_coefs[12][210] = 16'h0000;
	mel_filter_coefs[12][211] = 16'h0000;
	mel_filter_coefs[12][212] = 16'h0000;
	mel_filter_coefs[12][213] = 16'h0000;
	mel_filter_coefs[12][214] = 16'h0000;
	mel_filter_coefs[12][215] = 16'h0000;
	mel_filter_coefs[12][216] = 16'h0000;
	mel_filter_coefs[12][217] = 16'h0000;
	mel_filter_coefs[12][218] = 16'h0000;
	mel_filter_coefs[12][219] = 16'h0000;
	mel_filter_coefs[12][220] = 16'h0000;
	mel_filter_coefs[12][221] = 16'h0000;
	mel_filter_coefs[12][222] = 16'h0000;
	mel_filter_coefs[12][223] = 16'h0000;
	mel_filter_coefs[12][224] = 16'h0000;
	mel_filter_coefs[12][225] = 16'h0000;
	mel_filter_coefs[12][226] = 16'h0000;
	mel_filter_coefs[12][227] = 16'h0000;
	mel_filter_coefs[12][228] = 16'h0000;
	mel_filter_coefs[12][229] = 16'h0000;
	mel_filter_coefs[12][230] = 16'h0000;
	mel_filter_coefs[12][231] = 16'h0000;
	mel_filter_coefs[12][232] = 16'h0000;
	mel_filter_coefs[12][233] = 16'h0000;
	mel_filter_coefs[12][234] = 16'h0000;
	mel_filter_coefs[12][235] = 16'h0000;
	mel_filter_coefs[12][236] = 16'h0000;
	mel_filter_coefs[12][237] = 16'h0000;
	mel_filter_coefs[12][238] = 16'h0000;
	mel_filter_coefs[12][239] = 16'h0000;
	mel_filter_coefs[12][240] = 16'h0000;
	mel_filter_coefs[12][241] = 16'h0000;
	mel_filter_coefs[12][242] = 16'h0000;
	mel_filter_coefs[12][243] = 16'h0000;
	mel_filter_coefs[12][244] = 16'h0000;
	mel_filter_coefs[12][245] = 16'h0000;
	mel_filter_coefs[12][246] = 16'h0000;
	mel_filter_coefs[12][247] = 16'h0000;
	mel_filter_coefs[12][248] = 16'h0000;
	mel_filter_coefs[12][249] = 16'h0000;
	mel_filter_coefs[12][250] = 16'h0000;
	mel_filter_coefs[12][251] = 16'h0000;
	mel_filter_coefs[12][252] = 16'h0000;
	mel_filter_coefs[12][253] = 16'h0000;
	mel_filter_coefs[12][254] = 16'h0000;
	mel_filter_coefs[12][255] = 16'h0000;
	mel_filter_coefs[13][0] = 16'h0000;
	mel_filter_coefs[13][1] = 16'h0000;
	mel_filter_coefs[13][2] = 16'h0000;
	mel_filter_coefs[13][3] = 16'h0000;
	mel_filter_coefs[13][4] = 16'h0000;
	mel_filter_coefs[13][5] = 16'h0000;
	mel_filter_coefs[13][6] = 16'h0000;
	mel_filter_coefs[13][7] = 16'h0000;
	mel_filter_coefs[13][8] = 16'h0000;
	mel_filter_coefs[13][9] = 16'h0000;
	mel_filter_coefs[13][10] = 16'h0000;
	mel_filter_coefs[13][11] = 16'h0000;
	mel_filter_coefs[13][12] = 16'h0000;
	mel_filter_coefs[13][13] = 16'h0000;
	mel_filter_coefs[13][14] = 16'h0000;
	mel_filter_coefs[13][15] = 16'h0000;
	mel_filter_coefs[13][16] = 16'h0000;
	mel_filter_coefs[13][17] = 16'h0000;
	mel_filter_coefs[13][18] = 16'h0000;
	mel_filter_coefs[13][19] = 16'h0000;
	mel_filter_coefs[13][20] = 16'h0000;
	mel_filter_coefs[13][21] = 16'h0000;
	mel_filter_coefs[13][22] = 16'h0000;
	mel_filter_coefs[13][23] = 16'h0000;
	mel_filter_coefs[13][24] = 16'h0000;
	mel_filter_coefs[13][25] = 16'h0000;
	mel_filter_coefs[13][26] = 16'h0000;
	mel_filter_coefs[13][27] = 16'h0000;
	mel_filter_coefs[13][28] = 16'h1CA3;
	mel_filter_coefs[13][29] = 16'h4557;
	mel_filter_coefs[13][30] = 16'h6E0B;
	mel_filter_coefs[13][31] = 16'h6A9D;
	mel_filter_coefs[13][32] = 16'h4456;
	mel_filter_coefs[13][33] = 16'h1E0F;
	mel_filter_coefs[13][34] = 16'h0000;
	mel_filter_coefs[13][35] = 16'h0000;
	mel_filter_coefs[13][36] = 16'h0000;
	mel_filter_coefs[13][37] = 16'h0000;
	mel_filter_coefs[13][38] = 16'h0000;
	mel_filter_coefs[13][39] = 16'h0000;
	mel_filter_coefs[13][40] = 16'h0000;
	mel_filter_coefs[13][41] = 16'h0000;
	mel_filter_coefs[13][42] = 16'h0000;
	mel_filter_coefs[13][43] = 16'h0000;
	mel_filter_coefs[13][44] = 16'h0000;
	mel_filter_coefs[13][45] = 16'h0000;
	mel_filter_coefs[13][46] = 16'h0000;
	mel_filter_coefs[13][47] = 16'h0000;
	mel_filter_coefs[13][48] = 16'h0000;
	mel_filter_coefs[13][49] = 16'h0000;
	mel_filter_coefs[13][50] = 16'h0000;
	mel_filter_coefs[13][51] = 16'h0000;
	mel_filter_coefs[13][52] = 16'h0000;
	mel_filter_coefs[13][53] = 16'h0000;
	mel_filter_coefs[13][54] = 16'h0000;
	mel_filter_coefs[13][55] = 16'h0000;
	mel_filter_coefs[13][56] = 16'h0000;
	mel_filter_coefs[13][57] = 16'h0000;
	mel_filter_coefs[13][58] = 16'h0000;
	mel_filter_coefs[13][59] = 16'h0000;
	mel_filter_coefs[13][60] = 16'h0000;
	mel_filter_coefs[13][61] = 16'h0000;
	mel_filter_coefs[13][62] = 16'h0000;
	mel_filter_coefs[13][63] = 16'h0000;
	mel_filter_coefs[13][64] = 16'h0000;
	mel_filter_coefs[13][65] = 16'h0000;
	mel_filter_coefs[13][66] = 16'h0000;
	mel_filter_coefs[13][67] = 16'h0000;
	mel_filter_coefs[13][68] = 16'h0000;
	mel_filter_coefs[13][69] = 16'h0000;
	mel_filter_coefs[13][70] = 16'h0000;
	mel_filter_coefs[13][71] = 16'h0000;
	mel_filter_coefs[13][72] = 16'h0000;
	mel_filter_coefs[13][73] = 16'h0000;
	mel_filter_coefs[13][74] = 16'h0000;
	mel_filter_coefs[13][75] = 16'h0000;
	mel_filter_coefs[13][76] = 16'h0000;
	mel_filter_coefs[13][77] = 16'h0000;
	mel_filter_coefs[13][78] = 16'h0000;
	mel_filter_coefs[13][79] = 16'h0000;
	mel_filter_coefs[13][80] = 16'h0000;
	mel_filter_coefs[13][81] = 16'h0000;
	mel_filter_coefs[13][82] = 16'h0000;
	mel_filter_coefs[13][83] = 16'h0000;
	mel_filter_coefs[13][84] = 16'h0000;
	mel_filter_coefs[13][85] = 16'h0000;
	mel_filter_coefs[13][86] = 16'h0000;
	mel_filter_coefs[13][87] = 16'h0000;
	mel_filter_coefs[13][88] = 16'h0000;
	mel_filter_coefs[13][89] = 16'h0000;
	mel_filter_coefs[13][90] = 16'h0000;
	mel_filter_coefs[13][91] = 16'h0000;
	mel_filter_coefs[13][92] = 16'h0000;
	mel_filter_coefs[13][93] = 16'h0000;
	mel_filter_coefs[13][94] = 16'h0000;
	mel_filter_coefs[13][95] = 16'h0000;
	mel_filter_coefs[13][96] = 16'h0000;
	mel_filter_coefs[13][97] = 16'h0000;
	mel_filter_coefs[13][98] = 16'h0000;
	mel_filter_coefs[13][99] = 16'h0000;
	mel_filter_coefs[13][100] = 16'h0000;
	mel_filter_coefs[13][101] = 16'h0000;
	mel_filter_coefs[13][102] = 16'h0000;
	mel_filter_coefs[13][103] = 16'h0000;
	mel_filter_coefs[13][104] = 16'h0000;
	mel_filter_coefs[13][105] = 16'h0000;
	mel_filter_coefs[13][106] = 16'h0000;
	mel_filter_coefs[13][107] = 16'h0000;
	mel_filter_coefs[13][108] = 16'h0000;
	mel_filter_coefs[13][109] = 16'h0000;
	mel_filter_coefs[13][110] = 16'h0000;
	mel_filter_coefs[13][111] = 16'h0000;
	mel_filter_coefs[13][112] = 16'h0000;
	mel_filter_coefs[13][113] = 16'h0000;
	mel_filter_coefs[13][114] = 16'h0000;
	mel_filter_coefs[13][115] = 16'h0000;
	mel_filter_coefs[13][116] = 16'h0000;
	mel_filter_coefs[13][117] = 16'h0000;
	mel_filter_coefs[13][118] = 16'h0000;
	mel_filter_coefs[13][119] = 16'h0000;
	mel_filter_coefs[13][120] = 16'h0000;
	mel_filter_coefs[13][121] = 16'h0000;
	mel_filter_coefs[13][122] = 16'h0000;
	mel_filter_coefs[13][123] = 16'h0000;
	mel_filter_coefs[13][124] = 16'h0000;
	mel_filter_coefs[13][125] = 16'h0000;
	mel_filter_coefs[13][126] = 16'h0000;
	mel_filter_coefs[13][127] = 16'h0000;
	mel_filter_coefs[13][128] = 16'h0000;
	mel_filter_coefs[13][129] = 16'h0000;
	mel_filter_coefs[13][130] = 16'h0000;
	mel_filter_coefs[13][131] = 16'h0000;
	mel_filter_coefs[13][132] = 16'h0000;
	mel_filter_coefs[13][133] = 16'h0000;
	mel_filter_coefs[13][134] = 16'h0000;
	mel_filter_coefs[13][135] = 16'h0000;
	mel_filter_coefs[13][136] = 16'h0000;
	mel_filter_coefs[13][137] = 16'h0000;
	mel_filter_coefs[13][138] = 16'h0000;
	mel_filter_coefs[13][139] = 16'h0000;
	mel_filter_coefs[13][140] = 16'h0000;
	mel_filter_coefs[13][141] = 16'h0000;
	mel_filter_coefs[13][142] = 16'h0000;
	mel_filter_coefs[13][143] = 16'h0000;
	mel_filter_coefs[13][144] = 16'h0000;
	mel_filter_coefs[13][145] = 16'h0000;
	mel_filter_coefs[13][146] = 16'h0000;
	mel_filter_coefs[13][147] = 16'h0000;
	mel_filter_coefs[13][148] = 16'h0000;
	mel_filter_coefs[13][149] = 16'h0000;
	mel_filter_coefs[13][150] = 16'h0000;
	mel_filter_coefs[13][151] = 16'h0000;
	mel_filter_coefs[13][152] = 16'h0000;
	mel_filter_coefs[13][153] = 16'h0000;
	mel_filter_coefs[13][154] = 16'h0000;
	mel_filter_coefs[13][155] = 16'h0000;
	mel_filter_coefs[13][156] = 16'h0000;
	mel_filter_coefs[13][157] = 16'h0000;
	mel_filter_coefs[13][158] = 16'h0000;
	mel_filter_coefs[13][159] = 16'h0000;
	mel_filter_coefs[13][160] = 16'h0000;
	mel_filter_coefs[13][161] = 16'h0000;
	mel_filter_coefs[13][162] = 16'h0000;
	mel_filter_coefs[13][163] = 16'h0000;
	mel_filter_coefs[13][164] = 16'h0000;
	mel_filter_coefs[13][165] = 16'h0000;
	mel_filter_coefs[13][166] = 16'h0000;
	mel_filter_coefs[13][167] = 16'h0000;
	mel_filter_coefs[13][168] = 16'h0000;
	mel_filter_coefs[13][169] = 16'h0000;
	mel_filter_coefs[13][170] = 16'h0000;
	mel_filter_coefs[13][171] = 16'h0000;
	mel_filter_coefs[13][172] = 16'h0000;
	mel_filter_coefs[13][173] = 16'h0000;
	mel_filter_coefs[13][174] = 16'h0000;
	mel_filter_coefs[13][175] = 16'h0000;
	mel_filter_coefs[13][176] = 16'h0000;
	mel_filter_coefs[13][177] = 16'h0000;
	mel_filter_coefs[13][178] = 16'h0000;
	mel_filter_coefs[13][179] = 16'h0000;
	mel_filter_coefs[13][180] = 16'h0000;
	mel_filter_coefs[13][181] = 16'h0000;
	mel_filter_coefs[13][182] = 16'h0000;
	mel_filter_coefs[13][183] = 16'h0000;
	mel_filter_coefs[13][184] = 16'h0000;
	mel_filter_coefs[13][185] = 16'h0000;
	mel_filter_coefs[13][186] = 16'h0000;
	mel_filter_coefs[13][187] = 16'h0000;
	mel_filter_coefs[13][188] = 16'h0000;
	mel_filter_coefs[13][189] = 16'h0000;
	mel_filter_coefs[13][190] = 16'h0000;
	mel_filter_coefs[13][191] = 16'h0000;
	mel_filter_coefs[13][192] = 16'h0000;
	mel_filter_coefs[13][193] = 16'h0000;
	mel_filter_coefs[13][194] = 16'h0000;
	mel_filter_coefs[13][195] = 16'h0000;
	mel_filter_coefs[13][196] = 16'h0000;
	mel_filter_coefs[13][197] = 16'h0000;
	mel_filter_coefs[13][198] = 16'h0000;
	mel_filter_coefs[13][199] = 16'h0000;
	mel_filter_coefs[13][200] = 16'h0000;
	mel_filter_coefs[13][201] = 16'h0000;
	mel_filter_coefs[13][202] = 16'h0000;
	mel_filter_coefs[13][203] = 16'h0000;
	mel_filter_coefs[13][204] = 16'h0000;
	mel_filter_coefs[13][205] = 16'h0000;
	mel_filter_coefs[13][206] = 16'h0000;
	mel_filter_coefs[13][207] = 16'h0000;
	mel_filter_coefs[13][208] = 16'h0000;
	mel_filter_coefs[13][209] = 16'h0000;
	mel_filter_coefs[13][210] = 16'h0000;
	mel_filter_coefs[13][211] = 16'h0000;
	mel_filter_coefs[13][212] = 16'h0000;
	mel_filter_coefs[13][213] = 16'h0000;
	mel_filter_coefs[13][214] = 16'h0000;
	mel_filter_coefs[13][215] = 16'h0000;
	mel_filter_coefs[13][216] = 16'h0000;
	mel_filter_coefs[13][217] = 16'h0000;
	mel_filter_coefs[13][218] = 16'h0000;
	mel_filter_coefs[13][219] = 16'h0000;
	mel_filter_coefs[13][220] = 16'h0000;
	mel_filter_coefs[13][221] = 16'h0000;
	mel_filter_coefs[13][222] = 16'h0000;
	mel_filter_coefs[13][223] = 16'h0000;
	mel_filter_coefs[13][224] = 16'h0000;
	mel_filter_coefs[13][225] = 16'h0000;
	mel_filter_coefs[13][226] = 16'h0000;
	mel_filter_coefs[13][227] = 16'h0000;
	mel_filter_coefs[13][228] = 16'h0000;
	mel_filter_coefs[13][229] = 16'h0000;
	mel_filter_coefs[13][230] = 16'h0000;
	mel_filter_coefs[13][231] = 16'h0000;
	mel_filter_coefs[13][232] = 16'h0000;
	mel_filter_coefs[13][233] = 16'h0000;
	mel_filter_coefs[13][234] = 16'h0000;
	mel_filter_coefs[13][235] = 16'h0000;
	mel_filter_coefs[13][236] = 16'h0000;
	mel_filter_coefs[13][237] = 16'h0000;
	mel_filter_coefs[13][238] = 16'h0000;
	mel_filter_coefs[13][239] = 16'h0000;
	mel_filter_coefs[13][240] = 16'h0000;
	mel_filter_coefs[13][241] = 16'h0000;
	mel_filter_coefs[13][242] = 16'h0000;
	mel_filter_coefs[13][243] = 16'h0000;
	mel_filter_coefs[13][244] = 16'h0000;
	mel_filter_coefs[13][245] = 16'h0000;
	mel_filter_coefs[13][246] = 16'h0000;
	mel_filter_coefs[13][247] = 16'h0000;
	mel_filter_coefs[13][248] = 16'h0000;
	mel_filter_coefs[13][249] = 16'h0000;
	mel_filter_coefs[13][250] = 16'h0000;
	mel_filter_coefs[13][251] = 16'h0000;
	mel_filter_coefs[13][252] = 16'h0000;
	mel_filter_coefs[13][253] = 16'h0000;
	mel_filter_coefs[13][254] = 16'h0000;
	mel_filter_coefs[13][255] = 16'h0000;
	mel_filter_coefs[14][0] = 16'h0000;
	mel_filter_coefs[14][1] = 16'h0000;
	mel_filter_coefs[14][2] = 16'h0000;
	mel_filter_coefs[14][3] = 16'h0000;
	mel_filter_coefs[14][4] = 16'h0000;
	mel_filter_coefs[14][5] = 16'h0000;
	mel_filter_coefs[14][6] = 16'h0000;
	mel_filter_coefs[14][7] = 16'h0000;
	mel_filter_coefs[14][8] = 16'h0000;
	mel_filter_coefs[14][9] = 16'h0000;
	mel_filter_coefs[14][10] = 16'h0000;
	mel_filter_coefs[14][11] = 16'h0000;
	mel_filter_coefs[14][12] = 16'h0000;
	mel_filter_coefs[14][13] = 16'h0000;
	mel_filter_coefs[14][14] = 16'h0000;
	mel_filter_coefs[14][15] = 16'h0000;
	mel_filter_coefs[14][16] = 16'h0000;
	mel_filter_coefs[14][17] = 16'h0000;
	mel_filter_coefs[14][18] = 16'h0000;
	mel_filter_coefs[14][19] = 16'h0000;
	mel_filter_coefs[14][20] = 16'h0000;
	mel_filter_coefs[14][21] = 16'h0000;
	mel_filter_coefs[14][22] = 16'h0000;
	mel_filter_coefs[14][23] = 16'h0000;
	mel_filter_coefs[14][24] = 16'h0000;
	mel_filter_coefs[14][25] = 16'h0000;
	mel_filter_coefs[14][26] = 16'h0000;
	mel_filter_coefs[14][27] = 16'h0000;
	mel_filter_coefs[14][28] = 16'h0000;
	mel_filter_coefs[14][29] = 16'h0000;
	mel_filter_coefs[14][30] = 16'h0000;
	mel_filter_coefs[14][31] = 16'h1563;
	mel_filter_coefs[14][32] = 16'h3BAA;
	mel_filter_coefs[14][33] = 16'h61F1;
	mel_filter_coefs[14][34] = 16'h7846;
	mel_filter_coefs[14][35] = 16'h5448;
	mel_filter_coefs[14][36] = 16'h3049;
	mel_filter_coefs[14][37] = 16'h0C4B;
	mel_filter_coefs[14][38] = 16'h0000;
	mel_filter_coefs[14][39] = 16'h0000;
	mel_filter_coefs[14][40] = 16'h0000;
	mel_filter_coefs[14][41] = 16'h0000;
	mel_filter_coefs[14][42] = 16'h0000;
	mel_filter_coefs[14][43] = 16'h0000;
	mel_filter_coefs[14][44] = 16'h0000;
	mel_filter_coefs[14][45] = 16'h0000;
	mel_filter_coefs[14][46] = 16'h0000;
	mel_filter_coefs[14][47] = 16'h0000;
	mel_filter_coefs[14][48] = 16'h0000;
	mel_filter_coefs[14][49] = 16'h0000;
	mel_filter_coefs[14][50] = 16'h0000;
	mel_filter_coefs[14][51] = 16'h0000;
	mel_filter_coefs[14][52] = 16'h0000;
	mel_filter_coefs[14][53] = 16'h0000;
	mel_filter_coefs[14][54] = 16'h0000;
	mel_filter_coefs[14][55] = 16'h0000;
	mel_filter_coefs[14][56] = 16'h0000;
	mel_filter_coefs[14][57] = 16'h0000;
	mel_filter_coefs[14][58] = 16'h0000;
	mel_filter_coefs[14][59] = 16'h0000;
	mel_filter_coefs[14][60] = 16'h0000;
	mel_filter_coefs[14][61] = 16'h0000;
	mel_filter_coefs[14][62] = 16'h0000;
	mel_filter_coefs[14][63] = 16'h0000;
	mel_filter_coefs[14][64] = 16'h0000;
	mel_filter_coefs[14][65] = 16'h0000;
	mel_filter_coefs[14][66] = 16'h0000;
	mel_filter_coefs[14][67] = 16'h0000;
	mel_filter_coefs[14][68] = 16'h0000;
	mel_filter_coefs[14][69] = 16'h0000;
	mel_filter_coefs[14][70] = 16'h0000;
	mel_filter_coefs[14][71] = 16'h0000;
	mel_filter_coefs[14][72] = 16'h0000;
	mel_filter_coefs[14][73] = 16'h0000;
	mel_filter_coefs[14][74] = 16'h0000;
	mel_filter_coefs[14][75] = 16'h0000;
	mel_filter_coefs[14][76] = 16'h0000;
	mel_filter_coefs[14][77] = 16'h0000;
	mel_filter_coefs[14][78] = 16'h0000;
	mel_filter_coefs[14][79] = 16'h0000;
	mel_filter_coefs[14][80] = 16'h0000;
	mel_filter_coefs[14][81] = 16'h0000;
	mel_filter_coefs[14][82] = 16'h0000;
	mel_filter_coefs[14][83] = 16'h0000;
	mel_filter_coefs[14][84] = 16'h0000;
	mel_filter_coefs[14][85] = 16'h0000;
	mel_filter_coefs[14][86] = 16'h0000;
	mel_filter_coefs[14][87] = 16'h0000;
	mel_filter_coefs[14][88] = 16'h0000;
	mel_filter_coefs[14][89] = 16'h0000;
	mel_filter_coefs[14][90] = 16'h0000;
	mel_filter_coefs[14][91] = 16'h0000;
	mel_filter_coefs[14][92] = 16'h0000;
	mel_filter_coefs[14][93] = 16'h0000;
	mel_filter_coefs[14][94] = 16'h0000;
	mel_filter_coefs[14][95] = 16'h0000;
	mel_filter_coefs[14][96] = 16'h0000;
	mel_filter_coefs[14][97] = 16'h0000;
	mel_filter_coefs[14][98] = 16'h0000;
	mel_filter_coefs[14][99] = 16'h0000;
	mel_filter_coefs[14][100] = 16'h0000;
	mel_filter_coefs[14][101] = 16'h0000;
	mel_filter_coefs[14][102] = 16'h0000;
	mel_filter_coefs[14][103] = 16'h0000;
	mel_filter_coefs[14][104] = 16'h0000;
	mel_filter_coefs[14][105] = 16'h0000;
	mel_filter_coefs[14][106] = 16'h0000;
	mel_filter_coefs[14][107] = 16'h0000;
	mel_filter_coefs[14][108] = 16'h0000;
	mel_filter_coefs[14][109] = 16'h0000;
	mel_filter_coefs[14][110] = 16'h0000;
	mel_filter_coefs[14][111] = 16'h0000;
	mel_filter_coefs[14][112] = 16'h0000;
	mel_filter_coefs[14][113] = 16'h0000;
	mel_filter_coefs[14][114] = 16'h0000;
	mel_filter_coefs[14][115] = 16'h0000;
	mel_filter_coefs[14][116] = 16'h0000;
	mel_filter_coefs[14][117] = 16'h0000;
	mel_filter_coefs[14][118] = 16'h0000;
	mel_filter_coefs[14][119] = 16'h0000;
	mel_filter_coefs[14][120] = 16'h0000;
	mel_filter_coefs[14][121] = 16'h0000;
	mel_filter_coefs[14][122] = 16'h0000;
	mel_filter_coefs[14][123] = 16'h0000;
	mel_filter_coefs[14][124] = 16'h0000;
	mel_filter_coefs[14][125] = 16'h0000;
	mel_filter_coefs[14][126] = 16'h0000;
	mel_filter_coefs[14][127] = 16'h0000;
	mel_filter_coefs[14][128] = 16'h0000;
	mel_filter_coefs[14][129] = 16'h0000;
	mel_filter_coefs[14][130] = 16'h0000;
	mel_filter_coefs[14][131] = 16'h0000;
	mel_filter_coefs[14][132] = 16'h0000;
	mel_filter_coefs[14][133] = 16'h0000;
	mel_filter_coefs[14][134] = 16'h0000;
	mel_filter_coefs[14][135] = 16'h0000;
	mel_filter_coefs[14][136] = 16'h0000;
	mel_filter_coefs[14][137] = 16'h0000;
	mel_filter_coefs[14][138] = 16'h0000;
	mel_filter_coefs[14][139] = 16'h0000;
	mel_filter_coefs[14][140] = 16'h0000;
	mel_filter_coefs[14][141] = 16'h0000;
	mel_filter_coefs[14][142] = 16'h0000;
	mel_filter_coefs[14][143] = 16'h0000;
	mel_filter_coefs[14][144] = 16'h0000;
	mel_filter_coefs[14][145] = 16'h0000;
	mel_filter_coefs[14][146] = 16'h0000;
	mel_filter_coefs[14][147] = 16'h0000;
	mel_filter_coefs[14][148] = 16'h0000;
	mel_filter_coefs[14][149] = 16'h0000;
	mel_filter_coefs[14][150] = 16'h0000;
	mel_filter_coefs[14][151] = 16'h0000;
	mel_filter_coefs[14][152] = 16'h0000;
	mel_filter_coefs[14][153] = 16'h0000;
	mel_filter_coefs[14][154] = 16'h0000;
	mel_filter_coefs[14][155] = 16'h0000;
	mel_filter_coefs[14][156] = 16'h0000;
	mel_filter_coefs[14][157] = 16'h0000;
	mel_filter_coefs[14][158] = 16'h0000;
	mel_filter_coefs[14][159] = 16'h0000;
	mel_filter_coefs[14][160] = 16'h0000;
	mel_filter_coefs[14][161] = 16'h0000;
	mel_filter_coefs[14][162] = 16'h0000;
	mel_filter_coefs[14][163] = 16'h0000;
	mel_filter_coefs[14][164] = 16'h0000;
	mel_filter_coefs[14][165] = 16'h0000;
	mel_filter_coefs[14][166] = 16'h0000;
	mel_filter_coefs[14][167] = 16'h0000;
	mel_filter_coefs[14][168] = 16'h0000;
	mel_filter_coefs[14][169] = 16'h0000;
	mel_filter_coefs[14][170] = 16'h0000;
	mel_filter_coefs[14][171] = 16'h0000;
	mel_filter_coefs[14][172] = 16'h0000;
	mel_filter_coefs[14][173] = 16'h0000;
	mel_filter_coefs[14][174] = 16'h0000;
	mel_filter_coefs[14][175] = 16'h0000;
	mel_filter_coefs[14][176] = 16'h0000;
	mel_filter_coefs[14][177] = 16'h0000;
	mel_filter_coefs[14][178] = 16'h0000;
	mel_filter_coefs[14][179] = 16'h0000;
	mel_filter_coefs[14][180] = 16'h0000;
	mel_filter_coefs[14][181] = 16'h0000;
	mel_filter_coefs[14][182] = 16'h0000;
	mel_filter_coefs[14][183] = 16'h0000;
	mel_filter_coefs[14][184] = 16'h0000;
	mel_filter_coefs[14][185] = 16'h0000;
	mel_filter_coefs[14][186] = 16'h0000;
	mel_filter_coefs[14][187] = 16'h0000;
	mel_filter_coefs[14][188] = 16'h0000;
	mel_filter_coefs[14][189] = 16'h0000;
	mel_filter_coefs[14][190] = 16'h0000;
	mel_filter_coefs[14][191] = 16'h0000;
	mel_filter_coefs[14][192] = 16'h0000;
	mel_filter_coefs[14][193] = 16'h0000;
	mel_filter_coefs[14][194] = 16'h0000;
	mel_filter_coefs[14][195] = 16'h0000;
	mel_filter_coefs[14][196] = 16'h0000;
	mel_filter_coefs[14][197] = 16'h0000;
	mel_filter_coefs[14][198] = 16'h0000;
	mel_filter_coefs[14][199] = 16'h0000;
	mel_filter_coefs[14][200] = 16'h0000;
	mel_filter_coefs[14][201] = 16'h0000;
	mel_filter_coefs[14][202] = 16'h0000;
	mel_filter_coefs[14][203] = 16'h0000;
	mel_filter_coefs[14][204] = 16'h0000;
	mel_filter_coefs[14][205] = 16'h0000;
	mel_filter_coefs[14][206] = 16'h0000;
	mel_filter_coefs[14][207] = 16'h0000;
	mel_filter_coefs[14][208] = 16'h0000;
	mel_filter_coefs[14][209] = 16'h0000;
	mel_filter_coefs[14][210] = 16'h0000;
	mel_filter_coefs[14][211] = 16'h0000;
	mel_filter_coefs[14][212] = 16'h0000;
	mel_filter_coefs[14][213] = 16'h0000;
	mel_filter_coefs[14][214] = 16'h0000;
	mel_filter_coefs[14][215] = 16'h0000;
	mel_filter_coefs[14][216] = 16'h0000;
	mel_filter_coefs[14][217] = 16'h0000;
	mel_filter_coefs[14][218] = 16'h0000;
	mel_filter_coefs[14][219] = 16'h0000;
	mel_filter_coefs[14][220] = 16'h0000;
	mel_filter_coefs[14][221] = 16'h0000;
	mel_filter_coefs[14][222] = 16'h0000;
	mel_filter_coefs[14][223] = 16'h0000;
	mel_filter_coefs[14][224] = 16'h0000;
	mel_filter_coefs[14][225] = 16'h0000;
	mel_filter_coefs[14][226] = 16'h0000;
	mel_filter_coefs[14][227] = 16'h0000;
	mel_filter_coefs[14][228] = 16'h0000;
	mel_filter_coefs[14][229] = 16'h0000;
	mel_filter_coefs[14][230] = 16'h0000;
	mel_filter_coefs[14][231] = 16'h0000;
	mel_filter_coefs[14][232] = 16'h0000;
	mel_filter_coefs[14][233] = 16'h0000;
	mel_filter_coefs[14][234] = 16'h0000;
	mel_filter_coefs[14][235] = 16'h0000;
	mel_filter_coefs[14][236] = 16'h0000;
	mel_filter_coefs[14][237] = 16'h0000;
	mel_filter_coefs[14][238] = 16'h0000;
	mel_filter_coefs[14][239] = 16'h0000;
	mel_filter_coefs[14][240] = 16'h0000;
	mel_filter_coefs[14][241] = 16'h0000;
	mel_filter_coefs[14][242] = 16'h0000;
	mel_filter_coefs[14][243] = 16'h0000;
	mel_filter_coefs[14][244] = 16'h0000;
	mel_filter_coefs[14][245] = 16'h0000;
	mel_filter_coefs[14][246] = 16'h0000;
	mel_filter_coefs[14][247] = 16'h0000;
	mel_filter_coefs[14][248] = 16'h0000;
	mel_filter_coefs[14][249] = 16'h0000;
	mel_filter_coefs[14][250] = 16'h0000;
	mel_filter_coefs[14][251] = 16'h0000;
	mel_filter_coefs[14][252] = 16'h0000;
	mel_filter_coefs[14][253] = 16'h0000;
	mel_filter_coefs[14][254] = 16'h0000;
	mel_filter_coefs[14][255] = 16'h0000;
	mel_filter_coefs[15][0] = 16'h0000;
	mel_filter_coefs[15][1] = 16'h0000;
	mel_filter_coefs[15][2] = 16'h0000;
	mel_filter_coefs[15][3] = 16'h0000;
	mel_filter_coefs[15][4] = 16'h0000;
	mel_filter_coefs[15][5] = 16'h0000;
	mel_filter_coefs[15][6] = 16'h0000;
	mel_filter_coefs[15][7] = 16'h0000;
	mel_filter_coefs[15][8] = 16'h0000;
	mel_filter_coefs[15][9] = 16'h0000;
	mel_filter_coefs[15][10] = 16'h0000;
	mel_filter_coefs[15][11] = 16'h0000;
	mel_filter_coefs[15][12] = 16'h0000;
	mel_filter_coefs[15][13] = 16'h0000;
	mel_filter_coefs[15][14] = 16'h0000;
	mel_filter_coefs[15][15] = 16'h0000;
	mel_filter_coefs[15][16] = 16'h0000;
	mel_filter_coefs[15][17] = 16'h0000;
	mel_filter_coefs[15][18] = 16'h0000;
	mel_filter_coefs[15][19] = 16'h0000;
	mel_filter_coefs[15][20] = 16'h0000;
	mel_filter_coefs[15][21] = 16'h0000;
	mel_filter_coefs[15][22] = 16'h0000;
	mel_filter_coefs[15][23] = 16'h0000;
	mel_filter_coefs[15][24] = 16'h0000;
	mel_filter_coefs[15][25] = 16'h0000;
	mel_filter_coefs[15][26] = 16'h0000;
	mel_filter_coefs[15][27] = 16'h0000;
	mel_filter_coefs[15][28] = 16'h0000;
	mel_filter_coefs[15][29] = 16'h0000;
	mel_filter_coefs[15][30] = 16'h0000;
	mel_filter_coefs[15][31] = 16'h0000;
	mel_filter_coefs[15][32] = 16'h0000;
	mel_filter_coefs[15][33] = 16'h0000;
	mel_filter_coefs[15][34] = 16'h07BA;
	mel_filter_coefs[15][35] = 16'h2BB8;
	mel_filter_coefs[15][36] = 16'h4FB7;
	mel_filter_coefs[15][37] = 16'h73B5;
	mel_filter_coefs[15][38] = 16'h69B6;
	mel_filter_coefs[15][39] = 16'h47DD;
	mel_filter_coefs[15][40] = 16'h2603;
	mel_filter_coefs[15][41] = 16'h042A;
	mel_filter_coefs[15][42] = 16'h0000;
	mel_filter_coefs[15][43] = 16'h0000;
	mel_filter_coefs[15][44] = 16'h0000;
	mel_filter_coefs[15][45] = 16'h0000;
	mel_filter_coefs[15][46] = 16'h0000;
	mel_filter_coefs[15][47] = 16'h0000;
	mel_filter_coefs[15][48] = 16'h0000;
	mel_filter_coefs[15][49] = 16'h0000;
	mel_filter_coefs[15][50] = 16'h0000;
	mel_filter_coefs[15][51] = 16'h0000;
	mel_filter_coefs[15][52] = 16'h0000;
	mel_filter_coefs[15][53] = 16'h0000;
	mel_filter_coefs[15][54] = 16'h0000;
	mel_filter_coefs[15][55] = 16'h0000;
	mel_filter_coefs[15][56] = 16'h0000;
	mel_filter_coefs[15][57] = 16'h0000;
	mel_filter_coefs[15][58] = 16'h0000;
	mel_filter_coefs[15][59] = 16'h0000;
	mel_filter_coefs[15][60] = 16'h0000;
	mel_filter_coefs[15][61] = 16'h0000;
	mel_filter_coefs[15][62] = 16'h0000;
	mel_filter_coefs[15][63] = 16'h0000;
	mel_filter_coefs[15][64] = 16'h0000;
	mel_filter_coefs[15][65] = 16'h0000;
	mel_filter_coefs[15][66] = 16'h0000;
	mel_filter_coefs[15][67] = 16'h0000;
	mel_filter_coefs[15][68] = 16'h0000;
	mel_filter_coefs[15][69] = 16'h0000;
	mel_filter_coefs[15][70] = 16'h0000;
	mel_filter_coefs[15][71] = 16'h0000;
	mel_filter_coefs[15][72] = 16'h0000;
	mel_filter_coefs[15][73] = 16'h0000;
	mel_filter_coefs[15][74] = 16'h0000;
	mel_filter_coefs[15][75] = 16'h0000;
	mel_filter_coefs[15][76] = 16'h0000;
	mel_filter_coefs[15][77] = 16'h0000;
	mel_filter_coefs[15][78] = 16'h0000;
	mel_filter_coefs[15][79] = 16'h0000;
	mel_filter_coefs[15][80] = 16'h0000;
	mel_filter_coefs[15][81] = 16'h0000;
	mel_filter_coefs[15][82] = 16'h0000;
	mel_filter_coefs[15][83] = 16'h0000;
	mel_filter_coefs[15][84] = 16'h0000;
	mel_filter_coefs[15][85] = 16'h0000;
	mel_filter_coefs[15][86] = 16'h0000;
	mel_filter_coefs[15][87] = 16'h0000;
	mel_filter_coefs[15][88] = 16'h0000;
	mel_filter_coefs[15][89] = 16'h0000;
	mel_filter_coefs[15][90] = 16'h0000;
	mel_filter_coefs[15][91] = 16'h0000;
	mel_filter_coefs[15][92] = 16'h0000;
	mel_filter_coefs[15][93] = 16'h0000;
	mel_filter_coefs[15][94] = 16'h0000;
	mel_filter_coefs[15][95] = 16'h0000;
	mel_filter_coefs[15][96] = 16'h0000;
	mel_filter_coefs[15][97] = 16'h0000;
	mel_filter_coefs[15][98] = 16'h0000;
	mel_filter_coefs[15][99] = 16'h0000;
	mel_filter_coefs[15][100] = 16'h0000;
	mel_filter_coefs[15][101] = 16'h0000;
	mel_filter_coefs[15][102] = 16'h0000;
	mel_filter_coefs[15][103] = 16'h0000;
	mel_filter_coefs[15][104] = 16'h0000;
	mel_filter_coefs[15][105] = 16'h0000;
	mel_filter_coefs[15][106] = 16'h0000;
	mel_filter_coefs[15][107] = 16'h0000;
	mel_filter_coefs[15][108] = 16'h0000;
	mel_filter_coefs[15][109] = 16'h0000;
	mel_filter_coefs[15][110] = 16'h0000;
	mel_filter_coefs[15][111] = 16'h0000;
	mel_filter_coefs[15][112] = 16'h0000;
	mel_filter_coefs[15][113] = 16'h0000;
	mel_filter_coefs[15][114] = 16'h0000;
	mel_filter_coefs[15][115] = 16'h0000;
	mel_filter_coefs[15][116] = 16'h0000;
	mel_filter_coefs[15][117] = 16'h0000;
	mel_filter_coefs[15][118] = 16'h0000;
	mel_filter_coefs[15][119] = 16'h0000;
	mel_filter_coefs[15][120] = 16'h0000;
	mel_filter_coefs[15][121] = 16'h0000;
	mel_filter_coefs[15][122] = 16'h0000;
	mel_filter_coefs[15][123] = 16'h0000;
	mel_filter_coefs[15][124] = 16'h0000;
	mel_filter_coefs[15][125] = 16'h0000;
	mel_filter_coefs[15][126] = 16'h0000;
	mel_filter_coefs[15][127] = 16'h0000;
	mel_filter_coefs[15][128] = 16'h0000;
	mel_filter_coefs[15][129] = 16'h0000;
	mel_filter_coefs[15][130] = 16'h0000;
	mel_filter_coefs[15][131] = 16'h0000;
	mel_filter_coefs[15][132] = 16'h0000;
	mel_filter_coefs[15][133] = 16'h0000;
	mel_filter_coefs[15][134] = 16'h0000;
	mel_filter_coefs[15][135] = 16'h0000;
	mel_filter_coefs[15][136] = 16'h0000;
	mel_filter_coefs[15][137] = 16'h0000;
	mel_filter_coefs[15][138] = 16'h0000;
	mel_filter_coefs[15][139] = 16'h0000;
	mel_filter_coefs[15][140] = 16'h0000;
	mel_filter_coefs[15][141] = 16'h0000;
	mel_filter_coefs[15][142] = 16'h0000;
	mel_filter_coefs[15][143] = 16'h0000;
	mel_filter_coefs[15][144] = 16'h0000;
	mel_filter_coefs[15][145] = 16'h0000;
	mel_filter_coefs[15][146] = 16'h0000;
	mel_filter_coefs[15][147] = 16'h0000;
	mel_filter_coefs[15][148] = 16'h0000;
	mel_filter_coefs[15][149] = 16'h0000;
	mel_filter_coefs[15][150] = 16'h0000;
	mel_filter_coefs[15][151] = 16'h0000;
	mel_filter_coefs[15][152] = 16'h0000;
	mel_filter_coefs[15][153] = 16'h0000;
	mel_filter_coefs[15][154] = 16'h0000;
	mel_filter_coefs[15][155] = 16'h0000;
	mel_filter_coefs[15][156] = 16'h0000;
	mel_filter_coefs[15][157] = 16'h0000;
	mel_filter_coefs[15][158] = 16'h0000;
	mel_filter_coefs[15][159] = 16'h0000;
	mel_filter_coefs[15][160] = 16'h0000;
	mel_filter_coefs[15][161] = 16'h0000;
	mel_filter_coefs[15][162] = 16'h0000;
	mel_filter_coefs[15][163] = 16'h0000;
	mel_filter_coefs[15][164] = 16'h0000;
	mel_filter_coefs[15][165] = 16'h0000;
	mel_filter_coefs[15][166] = 16'h0000;
	mel_filter_coefs[15][167] = 16'h0000;
	mel_filter_coefs[15][168] = 16'h0000;
	mel_filter_coefs[15][169] = 16'h0000;
	mel_filter_coefs[15][170] = 16'h0000;
	mel_filter_coefs[15][171] = 16'h0000;
	mel_filter_coefs[15][172] = 16'h0000;
	mel_filter_coefs[15][173] = 16'h0000;
	mel_filter_coefs[15][174] = 16'h0000;
	mel_filter_coefs[15][175] = 16'h0000;
	mel_filter_coefs[15][176] = 16'h0000;
	mel_filter_coefs[15][177] = 16'h0000;
	mel_filter_coefs[15][178] = 16'h0000;
	mel_filter_coefs[15][179] = 16'h0000;
	mel_filter_coefs[15][180] = 16'h0000;
	mel_filter_coefs[15][181] = 16'h0000;
	mel_filter_coefs[15][182] = 16'h0000;
	mel_filter_coefs[15][183] = 16'h0000;
	mel_filter_coefs[15][184] = 16'h0000;
	mel_filter_coefs[15][185] = 16'h0000;
	mel_filter_coefs[15][186] = 16'h0000;
	mel_filter_coefs[15][187] = 16'h0000;
	mel_filter_coefs[15][188] = 16'h0000;
	mel_filter_coefs[15][189] = 16'h0000;
	mel_filter_coefs[15][190] = 16'h0000;
	mel_filter_coefs[15][191] = 16'h0000;
	mel_filter_coefs[15][192] = 16'h0000;
	mel_filter_coefs[15][193] = 16'h0000;
	mel_filter_coefs[15][194] = 16'h0000;
	mel_filter_coefs[15][195] = 16'h0000;
	mel_filter_coefs[15][196] = 16'h0000;
	mel_filter_coefs[15][197] = 16'h0000;
	mel_filter_coefs[15][198] = 16'h0000;
	mel_filter_coefs[15][199] = 16'h0000;
	mel_filter_coefs[15][200] = 16'h0000;
	mel_filter_coefs[15][201] = 16'h0000;
	mel_filter_coefs[15][202] = 16'h0000;
	mel_filter_coefs[15][203] = 16'h0000;
	mel_filter_coefs[15][204] = 16'h0000;
	mel_filter_coefs[15][205] = 16'h0000;
	mel_filter_coefs[15][206] = 16'h0000;
	mel_filter_coefs[15][207] = 16'h0000;
	mel_filter_coefs[15][208] = 16'h0000;
	mel_filter_coefs[15][209] = 16'h0000;
	mel_filter_coefs[15][210] = 16'h0000;
	mel_filter_coefs[15][211] = 16'h0000;
	mel_filter_coefs[15][212] = 16'h0000;
	mel_filter_coefs[15][213] = 16'h0000;
	mel_filter_coefs[15][214] = 16'h0000;
	mel_filter_coefs[15][215] = 16'h0000;
	mel_filter_coefs[15][216] = 16'h0000;
	mel_filter_coefs[15][217] = 16'h0000;
	mel_filter_coefs[15][218] = 16'h0000;
	mel_filter_coefs[15][219] = 16'h0000;
	mel_filter_coefs[15][220] = 16'h0000;
	mel_filter_coefs[15][221] = 16'h0000;
	mel_filter_coefs[15][222] = 16'h0000;
	mel_filter_coefs[15][223] = 16'h0000;
	mel_filter_coefs[15][224] = 16'h0000;
	mel_filter_coefs[15][225] = 16'h0000;
	mel_filter_coefs[15][226] = 16'h0000;
	mel_filter_coefs[15][227] = 16'h0000;
	mel_filter_coefs[15][228] = 16'h0000;
	mel_filter_coefs[15][229] = 16'h0000;
	mel_filter_coefs[15][230] = 16'h0000;
	mel_filter_coefs[15][231] = 16'h0000;
	mel_filter_coefs[15][232] = 16'h0000;
	mel_filter_coefs[15][233] = 16'h0000;
	mel_filter_coefs[15][234] = 16'h0000;
	mel_filter_coefs[15][235] = 16'h0000;
	mel_filter_coefs[15][236] = 16'h0000;
	mel_filter_coefs[15][237] = 16'h0000;
	mel_filter_coefs[15][238] = 16'h0000;
	mel_filter_coefs[15][239] = 16'h0000;
	mel_filter_coefs[15][240] = 16'h0000;
	mel_filter_coefs[15][241] = 16'h0000;
	mel_filter_coefs[15][242] = 16'h0000;
	mel_filter_coefs[15][243] = 16'h0000;
	mel_filter_coefs[15][244] = 16'h0000;
	mel_filter_coefs[15][245] = 16'h0000;
	mel_filter_coefs[15][246] = 16'h0000;
	mel_filter_coefs[15][247] = 16'h0000;
	mel_filter_coefs[15][248] = 16'h0000;
	mel_filter_coefs[15][249] = 16'h0000;
	mel_filter_coefs[15][250] = 16'h0000;
	mel_filter_coefs[15][251] = 16'h0000;
	mel_filter_coefs[15][252] = 16'h0000;
	mel_filter_coefs[15][253] = 16'h0000;
	mel_filter_coefs[15][254] = 16'h0000;
	mel_filter_coefs[15][255] = 16'h0000;
	mel_filter_coefs[16][0] = 16'h0000;
	mel_filter_coefs[16][1] = 16'h0000;
	mel_filter_coefs[16][2] = 16'h0000;
	mel_filter_coefs[16][3] = 16'h0000;
	mel_filter_coefs[16][4] = 16'h0000;
	mel_filter_coefs[16][5] = 16'h0000;
	mel_filter_coefs[16][6] = 16'h0000;
	mel_filter_coefs[16][7] = 16'h0000;
	mel_filter_coefs[16][8] = 16'h0000;
	mel_filter_coefs[16][9] = 16'h0000;
	mel_filter_coefs[16][10] = 16'h0000;
	mel_filter_coefs[16][11] = 16'h0000;
	mel_filter_coefs[16][12] = 16'h0000;
	mel_filter_coefs[16][13] = 16'h0000;
	mel_filter_coefs[16][14] = 16'h0000;
	mel_filter_coefs[16][15] = 16'h0000;
	mel_filter_coefs[16][16] = 16'h0000;
	mel_filter_coefs[16][17] = 16'h0000;
	mel_filter_coefs[16][18] = 16'h0000;
	mel_filter_coefs[16][19] = 16'h0000;
	mel_filter_coefs[16][20] = 16'h0000;
	mel_filter_coefs[16][21] = 16'h0000;
	mel_filter_coefs[16][22] = 16'h0000;
	mel_filter_coefs[16][23] = 16'h0000;
	mel_filter_coefs[16][24] = 16'h0000;
	mel_filter_coefs[16][25] = 16'h0000;
	mel_filter_coefs[16][26] = 16'h0000;
	mel_filter_coefs[16][27] = 16'h0000;
	mel_filter_coefs[16][28] = 16'h0000;
	mel_filter_coefs[16][29] = 16'h0000;
	mel_filter_coefs[16][30] = 16'h0000;
	mel_filter_coefs[16][31] = 16'h0000;
	mel_filter_coefs[16][32] = 16'h0000;
	mel_filter_coefs[16][33] = 16'h0000;
	mel_filter_coefs[16][34] = 16'h0000;
	mel_filter_coefs[16][35] = 16'h0000;
	mel_filter_coefs[16][36] = 16'h0000;
	mel_filter_coefs[16][37] = 16'h0000;
	mel_filter_coefs[16][38] = 16'h164A;
	mel_filter_coefs[16][39] = 16'h3823;
	mel_filter_coefs[16][40] = 16'h59FD;
	mel_filter_coefs[16][41] = 16'h7BD6;
	mel_filter_coefs[16][42] = 16'h6416;
	mel_filter_coefs[16][43] = 16'h4441;
	mel_filter_coefs[16][44] = 16'h246D;
	mel_filter_coefs[16][45] = 16'h0498;
	mel_filter_coefs[16][46] = 16'h0000;
	mel_filter_coefs[16][47] = 16'h0000;
	mel_filter_coefs[16][48] = 16'h0000;
	mel_filter_coefs[16][49] = 16'h0000;
	mel_filter_coefs[16][50] = 16'h0000;
	mel_filter_coefs[16][51] = 16'h0000;
	mel_filter_coefs[16][52] = 16'h0000;
	mel_filter_coefs[16][53] = 16'h0000;
	mel_filter_coefs[16][54] = 16'h0000;
	mel_filter_coefs[16][55] = 16'h0000;
	mel_filter_coefs[16][56] = 16'h0000;
	mel_filter_coefs[16][57] = 16'h0000;
	mel_filter_coefs[16][58] = 16'h0000;
	mel_filter_coefs[16][59] = 16'h0000;
	mel_filter_coefs[16][60] = 16'h0000;
	mel_filter_coefs[16][61] = 16'h0000;
	mel_filter_coefs[16][62] = 16'h0000;
	mel_filter_coefs[16][63] = 16'h0000;
	mel_filter_coefs[16][64] = 16'h0000;
	mel_filter_coefs[16][65] = 16'h0000;
	mel_filter_coefs[16][66] = 16'h0000;
	mel_filter_coefs[16][67] = 16'h0000;
	mel_filter_coefs[16][68] = 16'h0000;
	mel_filter_coefs[16][69] = 16'h0000;
	mel_filter_coefs[16][70] = 16'h0000;
	mel_filter_coefs[16][71] = 16'h0000;
	mel_filter_coefs[16][72] = 16'h0000;
	mel_filter_coefs[16][73] = 16'h0000;
	mel_filter_coefs[16][74] = 16'h0000;
	mel_filter_coefs[16][75] = 16'h0000;
	mel_filter_coefs[16][76] = 16'h0000;
	mel_filter_coefs[16][77] = 16'h0000;
	mel_filter_coefs[16][78] = 16'h0000;
	mel_filter_coefs[16][79] = 16'h0000;
	mel_filter_coefs[16][80] = 16'h0000;
	mel_filter_coefs[16][81] = 16'h0000;
	mel_filter_coefs[16][82] = 16'h0000;
	mel_filter_coefs[16][83] = 16'h0000;
	mel_filter_coefs[16][84] = 16'h0000;
	mel_filter_coefs[16][85] = 16'h0000;
	mel_filter_coefs[16][86] = 16'h0000;
	mel_filter_coefs[16][87] = 16'h0000;
	mel_filter_coefs[16][88] = 16'h0000;
	mel_filter_coefs[16][89] = 16'h0000;
	mel_filter_coefs[16][90] = 16'h0000;
	mel_filter_coefs[16][91] = 16'h0000;
	mel_filter_coefs[16][92] = 16'h0000;
	mel_filter_coefs[16][93] = 16'h0000;
	mel_filter_coefs[16][94] = 16'h0000;
	mel_filter_coefs[16][95] = 16'h0000;
	mel_filter_coefs[16][96] = 16'h0000;
	mel_filter_coefs[16][97] = 16'h0000;
	mel_filter_coefs[16][98] = 16'h0000;
	mel_filter_coefs[16][99] = 16'h0000;
	mel_filter_coefs[16][100] = 16'h0000;
	mel_filter_coefs[16][101] = 16'h0000;
	mel_filter_coefs[16][102] = 16'h0000;
	mel_filter_coefs[16][103] = 16'h0000;
	mel_filter_coefs[16][104] = 16'h0000;
	mel_filter_coefs[16][105] = 16'h0000;
	mel_filter_coefs[16][106] = 16'h0000;
	mel_filter_coefs[16][107] = 16'h0000;
	mel_filter_coefs[16][108] = 16'h0000;
	mel_filter_coefs[16][109] = 16'h0000;
	mel_filter_coefs[16][110] = 16'h0000;
	mel_filter_coefs[16][111] = 16'h0000;
	mel_filter_coefs[16][112] = 16'h0000;
	mel_filter_coefs[16][113] = 16'h0000;
	mel_filter_coefs[16][114] = 16'h0000;
	mel_filter_coefs[16][115] = 16'h0000;
	mel_filter_coefs[16][116] = 16'h0000;
	mel_filter_coefs[16][117] = 16'h0000;
	mel_filter_coefs[16][118] = 16'h0000;
	mel_filter_coefs[16][119] = 16'h0000;
	mel_filter_coefs[16][120] = 16'h0000;
	mel_filter_coefs[16][121] = 16'h0000;
	mel_filter_coefs[16][122] = 16'h0000;
	mel_filter_coefs[16][123] = 16'h0000;
	mel_filter_coefs[16][124] = 16'h0000;
	mel_filter_coefs[16][125] = 16'h0000;
	mel_filter_coefs[16][126] = 16'h0000;
	mel_filter_coefs[16][127] = 16'h0000;
	mel_filter_coefs[16][128] = 16'h0000;
	mel_filter_coefs[16][129] = 16'h0000;
	mel_filter_coefs[16][130] = 16'h0000;
	mel_filter_coefs[16][131] = 16'h0000;
	mel_filter_coefs[16][132] = 16'h0000;
	mel_filter_coefs[16][133] = 16'h0000;
	mel_filter_coefs[16][134] = 16'h0000;
	mel_filter_coefs[16][135] = 16'h0000;
	mel_filter_coefs[16][136] = 16'h0000;
	mel_filter_coefs[16][137] = 16'h0000;
	mel_filter_coefs[16][138] = 16'h0000;
	mel_filter_coefs[16][139] = 16'h0000;
	mel_filter_coefs[16][140] = 16'h0000;
	mel_filter_coefs[16][141] = 16'h0000;
	mel_filter_coefs[16][142] = 16'h0000;
	mel_filter_coefs[16][143] = 16'h0000;
	mel_filter_coefs[16][144] = 16'h0000;
	mel_filter_coefs[16][145] = 16'h0000;
	mel_filter_coefs[16][146] = 16'h0000;
	mel_filter_coefs[16][147] = 16'h0000;
	mel_filter_coefs[16][148] = 16'h0000;
	mel_filter_coefs[16][149] = 16'h0000;
	mel_filter_coefs[16][150] = 16'h0000;
	mel_filter_coefs[16][151] = 16'h0000;
	mel_filter_coefs[16][152] = 16'h0000;
	mel_filter_coefs[16][153] = 16'h0000;
	mel_filter_coefs[16][154] = 16'h0000;
	mel_filter_coefs[16][155] = 16'h0000;
	mel_filter_coefs[16][156] = 16'h0000;
	mel_filter_coefs[16][157] = 16'h0000;
	mel_filter_coefs[16][158] = 16'h0000;
	mel_filter_coefs[16][159] = 16'h0000;
	mel_filter_coefs[16][160] = 16'h0000;
	mel_filter_coefs[16][161] = 16'h0000;
	mel_filter_coefs[16][162] = 16'h0000;
	mel_filter_coefs[16][163] = 16'h0000;
	mel_filter_coefs[16][164] = 16'h0000;
	mel_filter_coefs[16][165] = 16'h0000;
	mel_filter_coefs[16][166] = 16'h0000;
	mel_filter_coefs[16][167] = 16'h0000;
	mel_filter_coefs[16][168] = 16'h0000;
	mel_filter_coefs[16][169] = 16'h0000;
	mel_filter_coefs[16][170] = 16'h0000;
	mel_filter_coefs[16][171] = 16'h0000;
	mel_filter_coefs[16][172] = 16'h0000;
	mel_filter_coefs[16][173] = 16'h0000;
	mel_filter_coefs[16][174] = 16'h0000;
	mel_filter_coefs[16][175] = 16'h0000;
	mel_filter_coefs[16][176] = 16'h0000;
	mel_filter_coefs[16][177] = 16'h0000;
	mel_filter_coefs[16][178] = 16'h0000;
	mel_filter_coefs[16][179] = 16'h0000;
	mel_filter_coefs[16][180] = 16'h0000;
	mel_filter_coefs[16][181] = 16'h0000;
	mel_filter_coefs[16][182] = 16'h0000;
	mel_filter_coefs[16][183] = 16'h0000;
	mel_filter_coefs[16][184] = 16'h0000;
	mel_filter_coefs[16][185] = 16'h0000;
	mel_filter_coefs[16][186] = 16'h0000;
	mel_filter_coefs[16][187] = 16'h0000;
	mel_filter_coefs[16][188] = 16'h0000;
	mel_filter_coefs[16][189] = 16'h0000;
	mel_filter_coefs[16][190] = 16'h0000;
	mel_filter_coefs[16][191] = 16'h0000;
	mel_filter_coefs[16][192] = 16'h0000;
	mel_filter_coefs[16][193] = 16'h0000;
	mel_filter_coefs[16][194] = 16'h0000;
	mel_filter_coefs[16][195] = 16'h0000;
	mel_filter_coefs[16][196] = 16'h0000;
	mel_filter_coefs[16][197] = 16'h0000;
	mel_filter_coefs[16][198] = 16'h0000;
	mel_filter_coefs[16][199] = 16'h0000;
	mel_filter_coefs[16][200] = 16'h0000;
	mel_filter_coefs[16][201] = 16'h0000;
	mel_filter_coefs[16][202] = 16'h0000;
	mel_filter_coefs[16][203] = 16'h0000;
	mel_filter_coefs[16][204] = 16'h0000;
	mel_filter_coefs[16][205] = 16'h0000;
	mel_filter_coefs[16][206] = 16'h0000;
	mel_filter_coefs[16][207] = 16'h0000;
	mel_filter_coefs[16][208] = 16'h0000;
	mel_filter_coefs[16][209] = 16'h0000;
	mel_filter_coefs[16][210] = 16'h0000;
	mel_filter_coefs[16][211] = 16'h0000;
	mel_filter_coefs[16][212] = 16'h0000;
	mel_filter_coefs[16][213] = 16'h0000;
	mel_filter_coefs[16][214] = 16'h0000;
	mel_filter_coefs[16][215] = 16'h0000;
	mel_filter_coefs[16][216] = 16'h0000;
	mel_filter_coefs[16][217] = 16'h0000;
	mel_filter_coefs[16][218] = 16'h0000;
	mel_filter_coefs[16][219] = 16'h0000;
	mel_filter_coefs[16][220] = 16'h0000;
	mel_filter_coefs[16][221] = 16'h0000;
	mel_filter_coefs[16][222] = 16'h0000;
	mel_filter_coefs[16][223] = 16'h0000;
	mel_filter_coefs[16][224] = 16'h0000;
	mel_filter_coefs[16][225] = 16'h0000;
	mel_filter_coefs[16][226] = 16'h0000;
	mel_filter_coefs[16][227] = 16'h0000;
	mel_filter_coefs[16][228] = 16'h0000;
	mel_filter_coefs[16][229] = 16'h0000;
	mel_filter_coefs[16][230] = 16'h0000;
	mel_filter_coefs[16][231] = 16'h0000;
	mel_filter_coefs[16][232] = 16'h0000;
	mel_filter_coefs[16][233] = 16'h0000;
	mel_filter_coefs[16][234] = 16'h0000;
	mel_filter_coefs[16][235] = 16'h0000;
	mel_filter_coefs[16][236] = 16'h0000;
	mel_filter_coefs[16][237] = 16'h0000;
	mel_filter_coefs[16][238] = 16'h0000;
	mel_filter_coefs[16][239] = 16'h0000;
	mel_filter_coefs[16][240] = 16'h0000;
	mel_filter_coefs[16][241] = 16'h0000;
	mel_filter_coefs[16][242] = 16'h0000;
	mel_filter_coefs[16][243] = 16'h0000;
	mel_filter_coefs[16][244] = 16'h0000;
	mel_filter_coefs[16][245] = 16'h0000;
	mel_filter_coefs[16][246] = 16'h0000;
	mel_filter_coefs[16][247] = 16'h0000;
	mel_filter_coefs[16][248] = 16'h0000;
	mel_filter_coefs[16][249] = 16'h0000;
	mel_filter_coefs[16][250] = 16'h0000;
	mel_filter_coefs[16][251] = 16'h0000;
	mel_filter_coefs[16][252] = 16'h0000;
	mel_filter_coefs[16][253] = 16'h0000;
	mel_filter_coefs[16][254] = 16'h0000;
	mel_filter_coefs[16][255] = 16'h0000;
	mel_filter_coefs[17][0] = 16'h0000;
	mel_filter_coefs[17][1] = 16'h0000;
	mel_filter_coefs[17][2] = 16'h0000;
	mel_filter_coefs[17][3] = 16'h0000;
	mel_filter_coefs[17][4] = 16'h0000;
	mel_filter_coefs[17][5] = 16'h0000;
	mel_filter_coefs[17][6] = 16'h0000;
	mel_filter_coefs[17][7] = 16'h0000;
	mel_filter_coefs[17][8] = 16'h0000;
	mel_filter_coefs[17][9] = 16'h0000;
	mel_filter_coefs[17][10] = 16'h0000;
	mel_filter_coefs[17][11] = 16'h0000;
	mel_filter_coefs[17][12] = 16'h0000;
	mel_filter_coefs[17][13] = 16'h0000;
	mel_filter_coefs[17][14] = 16'h0000;
	mel_filter_coefs[17][15] = 16'h0000;
	mel_filter_coefs[17][16] = 16'h0000;
	mel_filter_coefs[17][17] = 16'h0000;
	mel_filter_coefs[17][18] = 16'h0000;
	mel_filter_coefs[17][19] = 16'h0000;
	mel_filter_coefs[17][20] = 16'h0000;
	mel_filter_coefs[17][21] = 16'h0000;
	mel_filter_coefs[17][22] = 16'h0000;
	mel_filter_coefs[17][23] = 16'h0000;
	mel_filter_coefs[17][24] = 16'h0000;
	mel_filter_coefs[17][25] = 16'h0000;
	mel_filter_coefs[17][26] = 16'h0000;
	mel_filter_coefs[17][27] = 16'h0000;
	mel_filter_coefs[17][28] = 16'h0000;
	mel_filter_coefs[17][29] = 16'h0000;
	mel_filter_coefs[17][30] = 16'h0000;
	mel_filter_coefs[17][31] = 16'h0000;
	mel_filter_coefs[17][32] = 16'h0000;
	mel_filter_coefs[17][33] = 16'h0000;
	mel_filter_coefs[17][34] = 16'h0000;
	mel_filter_coefs[17][35] = 16'h0000;
	mel_filter_coefs[17][36] = 16'h0000;
	mel_filter_coefs[17][37] = 16'h0000;
	mel_filter_coefs[17][38] = 16'h0000;
	mel_filter_coefs[17][39] = 16'h0000;
	mel_filter_coefs[17][40] = 16'h0000;
	mel_filter_coefs[17][41] = 16'h0000;
	mel_filter_coefs[17][42] = 16'h1BEA;
	mel_filter_coefs[17][43] = 16'h3BBF;
	mel_filter_coefs[17][44] = 16'h5B93;
	mel_filter_coefs[17][45] = 16'h7B68;
	mel_filter_coefs[17][46] = 16'h6663;
	mel_filter_coefs[17][47] = 16'h4874;
	mel_filter_coefs[17][48] = 16'h2A85;
	mel_filter_coefs[17][49] = 16'h0C96;
	mel_filter_coefs[17][50] = 16'h0000;
	mel_filter_coefs[17][51] = 16'h0000;
	mel_filter_coefs[17][52] = 16'h0000;
	mel_filter_coefs[17][53] = 16'h0000;
	mel_filter_coefs[17][54] = 16'h0000;
	mel_filter_coefs[17][55] = 16'h0000;
	mel_filter_coefs[17][56] = 16'h0000;
	mel_filter_coefs[17][57] = 16'h0000;
	mel_filter_coefs[17][58] = 16'h0000;
	mel_filter_coefs[17][59] = 16'h0000;
	mel_filter_coefs[17][60] = 16'h0000;
	mel_filter_coefs[17][61] = 16'h0000;
	mel_filter_coefs[17][62] = 16'h0000;
	mel_filter_coefs[17][63] = 16'h0000;
	mel_filter_coefs[17][64] = 16'h0000;
	mel_filter_coefs[17][65] = 16'h0000;
	mel_filter_coefs[17][66] = 16'h0000;
	mel_filter_coefs[17][67] = 16'h0000;
	mel_filter_coefs[17][68] = 16'h0000;
	mel_filter_coefs[17][69] = 16'h0000;
	mel_filter_coefs[17][70] = 16'h0000;
	mel_filter_coefs[17][71] = 16'h0000;
	mel_filter_coefs[17][72] = 16'h0000;
	mel_filter_coefs[17][73] = 16'h0000;
	mel_filter_coefs[17][74] = 16'h0000;
	mel_filter_coefs[17][75] = 16'h0000;
	mel_filter_coefs[17][76] = 16'h0000;
	mel_filter_coefs[17][77] = 16'h0000;
	mel_filter_coefs[17][78] = 16'h0000;
	mel_filter_coefs[17][79] = 16'h0000;
	mel_filter_coefs[17][80] = 16'h0000;
	mel_filter_coefs[17][81] = 16'h0000;
	mel_filter_coefs[17][82] = 16'h0000;
	mel_filter_coefs[17][83] = 16'h0000;
	mel_filter_coefs[17][84] = 16'h0000;
	mel_filter_coefs[17][85] = 16'h0000;
	mel_filter_coefs[17][86] = 16'h0000;
	mel_filter_coefs[17][87] = 16'h0000;
	mel_filter_coefs[17][88] = 16'h0000;
	mel_filter_coefs[17][89] = 16'h0000;
	mel_filter_coefs[17][90] = 16'h0000;
	mel_filter_coefs[17][91] = 16'h0000;
	mel_filter_coefs[17][92] = 16'h0000;
	mel_filter_coefs[17][93] = 16'h0000;
	mel_filter_coefs[17][94] = 16'h0000;
	mel_filter_coefs[17][95] = 16'h0000;
	mel_filter_coefs[17][96] = 16'h0000;
	mel_filter_coefs[17][97] = 16'h0000;
	mel_filter_coefs[17][98] = 16'h0000;
	mel_filter_coefs[17][99] = 16'h0000;
	mel_filter_coefs[17][100] = 16'h0000;
	mel_filter_coefs[17][101] = 16'h0000;
	mel_filter_coefs[17][102] = 16'h0000;
	mel_filter_coefs[17][103] = 16'h0000;
	mel_filter_coefs[17][104] = 16'h0000;
	mel_filter_coefs[17][105] = 16'h0000;
	mel_filter_coefs[17][106] = 16'h0000;
	mel_filter_coefs[17][107] = 16'h0000;
	mel_filter_coefs[17][108] = 16'h0000;
	mel_filter_coefs[17][109] = 16'h0000;
	mel_filter_coefs[17][110] = 16'h0000;
	mel_filter_coefs[17][111] = 16'h0000;
	mel_filter_coefs[17][112] = 16'h0000;
	mel_filter_coefs[17][113] = 16'h0000;
	mel_filter_coefs[17][114] = 16'h0000;
	mel_filter_coefs[17][115] = 16'h0000;
	mel_filter_coefs[17][116] = 16'h0000;
	mel_filter_coefs[17][117] = 16'h0000;
	mel_filter_coefs[17][118] = 16'h0000;
	mel_filter_coefs[17][119] = 16'h0000;
	mel_filter_coefs[17][120] = 16'h0000;
	mel_filter_coefs[17][121] = 16'h0000;
	mel_filter_coefs[17][122] = 16'h0000;
	mel_filter_coefs[17][123] = 16'h0000;
	mel_filter_coefs[17][124] = 16'h0000;
	mel_filter_coefs[17][125] = 16'h0000;
	mel_filter_coefs[17][126] = 16'h0000;
	mel_filter_coefs[17][127] = 16'h0000;
	mel_filter_coefs[17][128] = 16'h0000;
	mel_filter_coefs[17][129] = 16'h0000;
	mel_filter_coefs[17][130] = 16'h0000;
	mel_filter_coefs[17][131] = 16'h0000;
	mel_filter_coefs[17][132] = 16'h0000;
	mel_filter_coefs[17][133] = 16'h0000;
	mel_filter_coefs[17][134] = 16'h0000;
	mel_filter_coefs[17][135] = 16'h0000;
	mel_filter_coefs[17][136] = 16'h0000;
	mel_filter_coefs[17][137] = 16'h0000;
	mel_filter_coefs[17][138] = 16'h0000;
	mel_filter_coefs[17][139] = 16'h0000;
	mel_filter_coefs[17][140] = 16'h0000;
	mel_filter_coefs[17][141] = 16'h0000;
	mel_filter_coefs[17][142] = 16'h0000;
	mel_filter_coefs[17][143] = 16'h0000;
	mel_filter_coefs[17][144] = 16'h0000;
	mel_filter_coefs[17][145] = 16'h0000;
	mel_filter_coefs[17][146] = 16'h0000;
	mel_filter_coefs[17][147] = 16'h0000;
	mel_filter_coefs[17][148] = 16'h0000;
	mel_filter_coefs[17][149] = 16'h0000;
	mel_filter_coefs[17][150] = 16'h0000;
	mel_filter_coefs[17][151] = 16'h0000;
	mel_filter_coefs[17][152] = 16'h0000;
	mel_filter_coefs[17][153] = 16'h0000;
	mel_filter_coefs[17][154] = 16'h0000;
	mel_filter_coefs[17][155] = 16'h0000;
	mel_filter_coefs[17][156] = 16'h0000;
	mel_filter_coefs[17][157] = 16'h0000;
	mel_filter_coefs[17][158] = 16'h0000;
	mel_filter_coefs[17][159] = 16'h0000;
	mel_filter_coefs[17][160] = 16'h0000;
	mel_filter_coefs[17][161] = 16'h0000;
	mel_filter_coefs[17][162] = 16'h0000;
	mel_filter_coefs[17][163] = 16'h0000;
	mel_filter_coefs[17][164] = 16'h0000;
	mel_filter_coefs[17][165] = 16'h0000;
	mel_filter_coefs[17][166] = 16'h0000;
	mel_filter_coefs[17][167] = 16'h0000;
	mel_filter_coefs[17][168] = 16'h0000;
	mel_filter_coefs[17][169] = 16'h0000;
	mel_filter_coefs[17][170] = 16'h0000;
	mel_filter_coefs[17][171] = 16'h0000;
	mel_filter_coefs[17][172] = 16'h0000;
	mel_filter_coefs[17][173] = 16'h0000;
	mel_filter_coefs[17][174] = 16'h0000;
	mel_filter_coefs[17][175] = 16'h0000;
	mel_filter_coefs[17][176] = 16'h0000;
	mel_filter_coefs[17][177] = 16'h0000;
	mel_filter_coefs[17][178] = 16'h0000;
	mel_filter_coefs[17][179] = 16'h0000;
	mel_filter_coefs[17][180] = 16'h0000;
	mel_filter_coefs[17][181] = 16'h0000;
	mel_filter_coefs[17][182] = 16'h0000;
	mel_filter_coefs[17][183] = 16'h0000;
	mel_filter_coefs[17][184] = 16'h0000;
	mel_filter_coefs[17][185] = 16'h0000;
	mel_filter_coefs[17][186] = 16'h0000;
	mel_filter_coefs[17][187] = 16'h0000;
	mel_filter_coefs[17][188] = 16'h0000;
	mel_filter_coefs[17][189] = 16'h0000;
	mel_filter_coefs[17][190] = 16'h0000;
	mel_filter_coefs[17][191] = 16'h0000;
	mel_filter_coefs[17][192] = 16'h0000;
	mel_filter_coefs[17][193] = 16'h0000;
	mel_filter_coefs[17][194] = 16'h0000;
	mel_filter_coefs[17][195] = 16'h0000;
	mel_filter_coefs[17][196] = 16'h0000;
	mel_filter_coefs[17][197] = 16'h0000;
	mel_filter_coefs[17][198] = 16'h0000;
	mel_filter_coefs[17][199] = 16'h0000;
	mel_filter_coefs[17][200] = 16'h0000;
	mel_filter_coefs[17][201] = 16'h0000;
	mel_filter_coefs[17][202] = 16'h0000;
	mel_filter_coefs[17][203] = 16'h0000;
	mel_filter_coefs[17][204] = 16'h0000;
	mel_filter_coefs[17][205] = 16'h0000;
	mel_filter_coefs[17][206] = 16'h0000;
	mel_filter_coefs[17][207] = 16'h0000;
	mel_filter_coefs[17][208] = 16'h0000;
	mel_filter_coefs[17][209] = 16'h0000;
	mel_filter_coefs[17][210] = 16'h0000;
	mel_filter_coefs[17][211] = 16'h0000;
	mel_filter_coefs[17][212] = 16'h0000;
	mel_filter_coefs[17][213] = 16'h0000;
	mel_filter_coefs[17][214] = 16'h0000;
	mel_filter_coefs[17][215] = 16'h0000;
	mel_filter_coefs[17][216] = 16'h0000;
	mel_filter_coefs[17][217] = 16'h0000;
	mel_filter_coefs[17][218] = 16'h0000;
	mel_filter_coefs[17][219] = 16'h0000;
	mel_filter_coefs[17][220] = 16'h0000;
	mel_filter_coefs[17][221] = 16'h0000;
	mel_filter_coefs[17][222] = 16'h0000;
	mel_filter_coefs[17][223] = 16'h0000;
	mel_filter_coefs[17][224] = 16'h0000;
	mel_filter_coefs[17][225] = 16'h0000;
	mel_filter_coefs[17][226] = 16'h0000;
	mel_filter_coefs[17][227] = 16'h0000;
	mel_filter_coefs[17][228] = 16'h0000;
	mel_filter_coefs[17][229] = 16'h0000;
	mel_filter_coefs[17][230] = 16'h0000;
	mel_filter_coefs[17][231] = 16'h0000;
	mel_filter_coefs[17][232] = 16'h0000;
	mel_filter_coefs[17][233] = 16'h0000;
	mel_filter_coefs[17][234] = 16'h0000;
	mel_filter_coefs[17][235] = 16'h0000;
	mel_filter_coefs[17][236] = 16'h0000;
	mel_filter_coefs[17][237] = 16'h0000;
	mel_filter_coefs[17][238] = 16'h0000;
	mel_filter_coefs[17][239] = 16'h0000;
	mel_filter_coefs[17][240] = 16'h0000;
	mel_filter_coefs[17][241] = 16'h0000;
	mel_filter_coefs[17][242] = 16'h0000;
	mel_filter_coefs[17][243] = 16'h0000;
	mel_filter_coefs[17][244] = 16'h0000;
	mel_filter_coefs[17][245] = 16'h0000;
	mel_filter_coefs[17][246] = 16'h0000;
	mel_filter_coefs[17][247] = 16'h0000;
	mel_filter_coefs[17][248] = 16'h0000;
	mel_filter_coefs[17][249] = 16'h0000;
	mel_filter_coefs[17][250] = 16'h0000;
	mel_filter_coefs[17][251] = 16'h0000;
	mel_filter_coefs[17][252] = 16'h0000;
	mel_filter_coefs[17][253] = 16'h0000;
	mel_filter_coefs[17][254] = 16'h0000;
	mel_filter_coefs[17][255] = 16'h0000;
	mel_filter_coefs[18][0] = 16'h0000;
	mel_filter_coefs[18][1] = 16'h0000;
	mel_filter_coefs[18][2] = 16'h0000;
	mel_filter_coefs[18][3] = 16'h0000;
	mel_filter_coefs[18][4] = 16'h0000;
	mel_filter_coefs[18][5] = 16'h0000;
	mel_filter_coefs[18][6] = 16'h0000;
	mel_filter_coefs[18][7] = 16'h0000;
	mel_filter_coefs[18][8] = 16'h0000;
	mel_filter_coefs[18][9] = 16'h0000;
	mel_filter_coefs[18][10] = 16'h0000;
	mel_filter_coefs[18][11] = 16'h0000;
	mel_filter_coefs[18][12] = 16'h0000;
	mel_filter_coefs[18][13] = 16'h0000;
	mel_filter_coefs[18][14] = 16'h0000;
	mel_filter_coefs[18][15] = 16'h0000;
	mel_filter_coefs[18][16] = 16'h0000;
	mel_filter_coefs[18][17] = 16'h0000;
	mel_filter_coefs[18][18] = 16'h0000;
	mel_filter_coefs[18][19] = 16'h0000;
	mel_filter_coefs[18][20] = 16'h0000;
	mel_filter_coefs[18][21] = 16'h0000;
	mel_filter_coefs[18][22] = 16'h0000;
	mel_filter_coefs[18][23] = 16'h0000;
	mel_filter_coefs[18][24] = 16'h0000;
	mel_filter_coefs[18][25] = 16'h0000;
	mel_filter_coefs[18][26] = 16'h0000;
	mel_filter_coefs[18][27] = 16'h0000;
	mel_filter_coefs[18][28] = 16'h0000;
	mel_filter_coefs[18][29] = 16'h0000;
	mel_filter_coefs[18][30] = 16'h0000;
	mel_filter_coefs[18][31] = 16'h0000;
	mel_filter_coefs[18][32] = 16'h0000;
	mel_filter_coefs[18][33] = 16'h0000;
	mel_filter_coefs[18][34] = 16'h0000;
	mel_filter_coefs[18][35] = 16'h0000;
	mel_filter_coefs[18][36] = 16'h0000;
	mel_filter_coefs[18][37] = 16'h0000;
	mel_filter_coefs[18][38] = 16'h0000;
	mel_filter_coefs[18][39] = 16'h0000;
	mel_filter_coefs[18][40] = 16'h0000;
	mel_filter_coefs[18][41] = 16'h0000;
	mel_filter_coefs[18][42] = 16'h0000;
	mel_filter_coefs[18][43] = 16'h0000;
	mel_filter_coefs[18][44] = 16'h0000;
	mel_filter_coefs[18][45] = 16'h0000;
	mel_filter_coefs[18][46] = 16'h199D;
	mel_filter_coefs[18][47] = 16'h378C;
	mel_filter_coefs[18][48] = 16'h557B;
	mel_filter_coefs[18][49] = 16'h736A;
	mel_filter_coefs[18][50] = 16'h6FB0;
	mel_filter_coefs[18][51] = 16'h538A;
	mel_filter_coefs[18][52] = 16'h3764;
	mel_filter_coefs[18][53] = 16'h1B3E;
	mel_filter_coefs[18][54] = 16'h0000;
	mel_filter_coefs[18][55] = 16'h0000;
	mel_filter_coefs[18][56] = 16'h0000;
	mel_filter_coefs[18][57] = 16'h0000;
	mel_filter_coefs[18][58] = 16'h0000;
	mel_filter_coefs[18][59] = 16'h0000;
	mel_filter_coefs[18][60] = 16'h0000;
	mel_filter_coefs[18][61] = 16'h0000;
	mel_filter_coefs[18][62] = 16'h0000;
	mel_filter_coefs[18][63] = 16'h0000;
	mel_filter_coefs[18][64] = 16'h0000;
	mel_filter_coefs[18][65] = 16'h0000;
	mel_filter_coefs[18][66] = 16'h0000;
	mel_filter_coefs[18][67] = 16'h0000;
	mel_filter_coefs[18][68] = 16'h0000;
	mel_filter_coefs[18][69] = 16'h0000;
	mel_filter_coefs[18][70] = 16'h0000;
	mel_filter_coefs[18][71] = 16'h0000;
	mel_filter_coefs[18][72] = 16'h0000;
	mel_filter_coefs[18][73] = 16'h0000;
	mel_filter_coefs[18][74] = 16'h0000;
	mel_filter_coefs[18][75] = 16'h0000;
	mel_filter_coefs[18][76] = 16'h0000;
	mel_filter_coefs[18][77] = 16'h0000;
	mel_filter_coefs[18][78] = 16'h0000;
	mel_filter_coefs[18][79] = 16'h0000;
	mel_filter_coefs[18][80] = 16'h0000;
	mel_filter_coefs[18][81] = 16'h0000;
	mel_filter_coefs[18][82] = 16'h0000;
	mel_filter_coefs[18][83] = 16'h0000;
	mel_filter_coefs[18][84] = 16'h0000;
	mel_filter_coefs[18][85] = 16'h0000;
	mel_filter_coefs[18][86] = 16'h0000;
	mel_filter_coefs[18][87] = 16'h0000;
	mel_filter_coefs[18][88] = 16'h0000;
	mel_filter_coefs[18][89] = 16'h0000;
	mel_filter_coefs[18][90] = 16'h0000;
	mel_filter_coefs[18][91] = 16'h0000;
	mel_filter_coefs[18][92] = 16'h0000;
	mel_filter_coefs[18][93] = 16'h0000;
	mel_filter_coefs[18][94] = 16'h0000;
	mel_filter_coefs[18][95] = 16'h0000;
	mel_filter_coefs[18][96] = 16'h0000;
	mel_filter_coefs[18][97] = 16'h0000;
	mel_filter_coefs[18][98] = 16'h0000;
	mel_filter_coefs[18][99] = 16'h0000;
	mel_filter_coefs[18][100] = 16'h0000;
	mel_filter_coefs[18][101] = 16'h0000;
	mel_filter_coefs[18][102] = 16'h0000;
	mel_filter_coefs[18][103] = 16'h0000;
	mel_filter_coefs[18][104] = 16'h0000;
	mel_filter_coefs[18][105] = 16'h0000;
	mel_filter_coefs[18][106] = 16'h0000;
	mel_filter_coefs[18][107] = 16'h0000;
	mel_filter_coefs[18][108] = 16'h0000;
	mel_filter_coefs[18][109] = 16'h0000;
	mel_filter_coefs[18][110] = 16'h0000;
	mel_filter_coefs[18][111] = 16'h0000;
	mel_filter_coefs[18][112] = 16'h0000;
	mel_filter_coefs[18][113] = 16'h0000;
	mel_filter_coefs[18][114] = 16'h0000;
	mel_filter_coefs[18][115] = 16'h0000;
	mel_filter_coefs[18][116] = 16'h0000;
	mel_filter_coefs[18][117] = 16'h0000;
	mel_filter_coefs[18][118] = 16'h0000;
	mel_filter_coefs[18][119] = 16'h0000;
	mel_filter_coefs[18][120] = 16'h0000;
	mel_filter_coefs[18][121] = 16'h0000;
	mel_filter_coefs[18][122] = 16'h0000;
	mel_filter_coefs[18][123] = 16'h0000;
	mel_filter_coefs[18][124] = 16'h0000;
	mel_filter_coefs[18][125] = 16'h0000;
	mel_filter_coefs[18][126] = 16'h0000;
	mel_filter_coefs[18][127] = 16'h0000;
	mel_filter_coefs[18][128] = 16'h0000;
	mel_filter_coefs[18][129] = 16'h0000;
	mel_filter_coefs[18][130] = 16'h0000;
	mel_filter_coefs[18][131] = 16'h0000;
	mel_filter_coefs[18][132] = 16'h0000;
	mel_filter_coefs[18][133] = 16'h0000;
	mel_filter_coefs[18][134] = 16'h0000;
	mel_filter_coefs[18][135] = 16'h0000;
	mel_filter_coefs[18][136] = 16'h0000;
	mel_filter_coefs[18][137] = 16'h0000;
	mel_filter_coefs[18][138] = 16'h0000;
	mel_filter_coefs[18][139] = 16'h0000;
	mel_filter_coefs[18][140] = 16'h0000;
	mel_filter_coefs[18][141] = 16'h0000;
	mel_filter_coefs[18][142] = 16'h0000;
	mel_filter_coefs[18][143] = 16'h0000;
	mel_filter_coefs[18][144] = 16'h0000;
	mel_filter_coefs[18][145] = 16'h0000;
	mel_filter_coefs[18][146] = 16'h0000;
	mel_filter_coefs[18][147] = 16'h0000;
	mel_filter_coefs[18][148] = 16'h0000;
	mel_filter_coefs[18][149] = 16'h0000;
	mel_filter_coefs[18][150] = 16'h0000;
	mel_filter_coefs[18][151] = 16'h0000;
	mel_filter_coefs[18][152] = 16'h0000;
	mel_filter_coefs[18][153] = 16'h0000;
	mel_filter_coefs[18][154] = 16'h0000;
	mel_filter_coefs[18][155] = 16'h0000;
	mel_filter_coefs[18][156] = 16'h0000;
	mel_filter_coefs[18][157] = 16'h0000;
	mel_filter_coefs[18][158] = 16'h0000;
	mel_filter_coefs[18][159] = 16'h0000;
	mel_filter_coefs[18][160] = 16'h0000;
	mel_filter_coefs[18][161] = 16'h0000;
	mel_filter_coefs[18][162] = 16'h0000;
	mel_filter_coefs[18][163] = 16'h0000;
	mel_filter_coefs[18][164] = 16'h0000;
	mel_filter_coefs[18][165] = 16'h0000;
	mel_filter_coefs[18][166] = 16'h0000;
	mel_filter_coefs[18][167] = 16'h0000;
	mel_filter_coefs[18][168] = 16'h0000;
	mel_filter_coefs[18][169] = 16'h0000;
	mel_filter_coefs[18][170] = 16'h0000;
	mel_filter_coefs[18][171] = 16'h0000;
	mel_filter_coefs[18][172] = 16'h0000;
	mel_filter_coefs[18][173] = 16'h0000;
	mel_filter_coefs[18][174] = 16'h0000;
	mel_filter_coefs[18][175] = 16'h0000;
	mel_filter_coefs[18][176] = 16'h0000;
	mel_filter_coefs[18][177] = 16'h0000;
	mel_filter_coefs[18][178] = 16'h0000;
	mel_filter_coefs[18][179] = 16'h0000;
	mel_filter_coefs[18][180] = 16'h0000;
	mel_filter_coefs[18][181] = 16'h0000;
	mel_filter_coefs[18][182] = 16'h0000;
	mel_filter_coefs[18][183] = 16'h0000;
	mel_filter_coefs[18][184] = 16'h0000;
	mel_filter_coefs[18][185] = 16'h0000;
	mel_filter_coefs[18][186] = 16'h0000;
	mel_filter_coefs[18][187] = 16'h0000;
	mel_filter_coefs[18][188] = 16'h0000;
	mel_filter_coefs[18][189] = 16'h0000;
	mel_filter_coefs[18][190] = 16'h0000;
	mel_filter_coefs[18][191] = 16'h0000;
	mel_filter_coefs[18][192] = 16'h0000;
	mel_filter_coefs[18][193] = 16'h0000;
	mel_filter_coefs[18][194] = 16'h0000;
	mel_filter_coefs[18][195] = 16'h0000;
	mel_filter_coefs[18][196] = 16'h0000;
	mel_filter_coefs[18][197] = 16'h0000;
	mel_filter_coefs[18][198] = 16'h0000;
	mel_filter_coefs[18][199] = 16'h0000;
	mel_filter_coefs[18][200] = 16'h0000;
	mel_filter_coefs[18][201] = 16'h0000;
	mel_filter_coefs[18][202] = 16'h0000;
	mel_filter_coefs[18][203] = 16'h0000;
	mel_filter_coefs[18][204] = 16'h0000;
	mel_filter_coefs[18][205] = 16'h0000;
	mel_filter_coefs[18][206] = 16'h0000;
	mel_filter_coefs[18][207] = 16'h0000;
	mel_filter_coefs[18][208] = 16'h0000;
	mel_filter_coefs[18][209] = 16'h0000;
	mel_filter_coefs[18][210] = 16'h0000;
	mel_filter_coefs[18][211] = 16'h0000;
	mel_filter_coefs[18][212] = 16'h0000;
	mel_filter_coefs[18][213] = 16'h0000;
	mel_filter_coefs[18][214] = 16'h0000;
	mel_filter_coefs[18][215] = 16'h0000;
	mel_filter_coefs[18][216] = 16'h0000;
	mel_filter_coefs[18][217] = 16'h0000;
	mel_filter_coefs[18][218] = 16'h0000;
	mel_filter_coefs[18][219] = 16'h0000;
	mel_filter_coefs[18][220] = 16'h0000;
	mel_filter_coefs[18][221] = 16'h0000;
	mel_filter_coefs[18][222] = 16'h0000;
	mel_filter_coefs[18][223] = 16'h0000;
	mel_filter_coefs[18][224] = 16'h0000;
	mel_filter_coefs[18][225] = 16'h0000;
	mel_filter_coefs[18][226] = 16'h0000;
	mel_filter_coefs[18][227] = 16'h0000;
	mel_filter_coefs[18][228] = 16'h0000;
	mel_filter_coefs[18][229] = 16'h0000;
	mel_filter_coefs[18][230] = 16'h0000;
	mel_filter_coefs[18][231] = 16'h0000;
	mel_filter_coefs[18][232] = 16'h0000;
	mel_filter_coefs[18][233] = 16'h0000;
	mel_filter_coefs[18][234] = 16'h0000;
	mel_filter_coefs[18][235] = 16'h0000;
	mel_filter_coefs[18][236] = 16'h0000;
	mel_filter_coefs[18][237] = 16'h0000;
	mel_filter_coefs[18][238] = 16'h0000;
	mel_filter_coefs[18][239] = 16'h0000;
	mel_filter_coefs[18][240] = 16'h0000;
	mel_filter_coefs[18][241] = 16'h0000;
	mel_filter_coefs[18][242] = 16'h0000;
	mel_filter_coefs[18][243] = 16'h0000;
	mel_filter_coefs[18][244] = 16'h0000;
	mel_filter_coefs[18][245] = 16'h0000;
	mel_filter_coefs[18][246] = 16'h0000;
	mel_filter_coefs[18][247] = 16'h0000;
	mel_filter_coefs[18][248] = 16'h0000;
	mel_filter_coefs[18][249] = 16'h0000;
	mel_filter_coefs[18][250] = 16'h0000;
	mel_filter_coefs[18][251] = 16'h0000;
	mel_filter_coefs[18][252] = 16'h0000;
	mel_filter_coefs[18][253] = 16'h0000;
	mel_filter_coefs[18][254] = 16'h0000;
	mel_filter_coefs[18][255] = 16'h0000;
	mel_filter_coefs[19][0] = 16'h0000;
	mel_filter_coefs[19][1] = 16'h0000;
	mel_filter_coefs[19][2] = 16'h0000;
	mel_filter_coefs[19][3] = 16'h0000;
	mel_filter_coefs[19][4] = 16'h0000;
	mel_filter_coefs[19][5] = 16'h0000;
	mel_filter_coefs[19][6] = 16'h0000;
	mel_filter_coefs[19][7] = 16'h0000;
	mel_filter_coefs[19][8] = 16'h0000;
	mel_filter_coefs[19][9] = 16'h0000;
	mel_filter_coefs[19][10] = 16'h0000;
	mel_filter_coefs[19][11] = 16'h0000;
	mel_filter_coefs[19][12] = 16'h0000;
	mel_filter_coefs[19][13] = 16'h0000;
	mel_filter_coefs[19][14] = 16'h0000;
	mel_filter_coefs[19][15] = 16'h0000;
	mel_filter_coefs[19][16] = 16'h0000;
	mel_filter_coefs[19][17] = 16'h0000;
	mel_filter_coefs[19][18] = 16'h0000;
	mel_filter_coefs[19][19] = 16'h0000;
	mel_filter_coefs[19][20] = 16'h0000;
	mel_filter_coefs[19][21] = 16'h0000;
	mel_filter_coefs[19][22] = 16'h0000;
	mel_filter_coefs[19][23] = 16'h0000;
	mel_filter_coefs[19][24] = 16'h0000;
	mel_filter_coefs[19][25] = 16'h0000;
	mel_filter_coefs[19][26] = 16'h0000;
	mel_filter_coefs[19][27] = 16'h0000;
	mel_filter_coefs[19][28] = 16'h0000;
	mel_filter_coefs[19][29] = 16'h0000;
	mel_filter_coefs[19][30] = 16'h0000;
	mel_filter_coefs[19][31] = 16'h0000;
	mel_filter_coefs[19][32] = 16'h0000;
	mel_filter_coefs[19][33] = 16'h0000;
	mel_filter_coefs[19][34] = 16'h0000;
	mel_filter_coefs[19][35] = 16'h0000;
	mel_filter_coefs[19][36] = 16'h0000;
	mel_filter_coefs[19][37] = 16'h0000;
	mel_filter_coefs[19][38] = 16'h0000;
	mel_filter_coefs[19][39] = 16'h0000;
	mel_filter_coefs[19][40] = 16'h0000;
	mel_filter_coefs[19][41] = 16'h0000;
	mel_filter_coefs[19][42] = 16'h0000;
	mel_filter_coefs[19][43] = 16'h0000;
	mel_filter_coefs[19][44] = 16'h0000;
	mel_filter_coefs[19][45] = 16'h0000;
	mel_filter_coefs[19][46] = 16'h0000;
	mel_filter_coefs[19][47] = 16'h0000;
	mel_filter_coefs[19][48] = 16'h0000;
	mel_filter_coefs[19][49] = 16'h0000;
	mel_filter_coefs[19][50] = 16'h1050;
	mel_filter_coefs[19][51] = 16'h2C76;
	mel_filter_coefs[19][52] = 16'h489C;
	mel_filter_coefs[19][53] = 16'h64C2;
	mel_filter_coefs[19][54] = 16'h7F26;
	mel_filter_coefs[19][55] = 16'h64AD;
	mel_filter_coefs[19][56] = 16'h4A35;
	mel_filter_coefs[19][57] = 16'h2FBC;
	mel_filter_coefs[19][58] = 16'h1544;
	mel_filter_coefs[19][59] = 16'h0000;
	mel_filter_coefs[19][60] = 16'h0000;
	mel_filter_coefs[19][61] = 16'h0000;
	mel_filter_coefs[19][62] = 16'h0000;
	mel_filter_coefs[19][63] = 16'h0000;
	mel_filter_coefs[19][64] = 16'h0000;
	mel_filter_coefs[19][65] = 16'h0000;
	mel_filter_coefs[19][66] = 16'h0000;
	mel_filter_coefs[19][67] = 16'h0000;
	mel_filter_coefs[19][68] = 16'h0000;
	mel_filter_coefs[19][69] = 16'h0000;
	mel_filter_coefs[19][70] = 16'h0000;
	mel_filter_coefs[19][71] = 16'h0000;
	mel_filter_coefs[19][72] = 16'h0000;
	mel_filter_coefs[19][73] = 16'h0000;
	mel_filter_coefs[19][74] = 16'h0000;
	mel_filter_coefs[19][75] = 16'h0000;
	mel_filter_coefs[19][76] = 16'h0000;
	mel_filter_coefs[19][77] = 16'h0000;
	mel_filter_coefs[19][78] = 16'h0000;
	mel_filter_coefs[19][79] = 16'h0000;
	mel_filter_coefs[19][80] = 16'h0000;
	mel_filter_coefs[19][81] = 16'h0000;
	mel_filter_coefs[19][82] = 16'h0000;
	mel_filter_coefs[19][83] = 16'h0000;
	mel_filter_coefs[19][84] = 16'h0000;
	mel_filter_coefs[19][85] = 16'h0000;
	mel_filter_coefs[19][86] = 16'h0000;
	mel_filter_coefs[19][87] = 16'h0000;
	mel_filter_coefs[19][88] = 16'h0000;
	mel_filter_coefs[19][89] = 16'h0000;
	mel_filter_coefs[19][90] = 16'h0000;
	mel_filter_coefs[19][91] = 16'h0000;
	mel_filter_coefs[19][92] = 16'h0000;
	mel_filter_coefs[19][93] = 16'h0000;
	mel_filter_coefs[19][94] = 16'h0000;
	mel_filter_coefs[19][95] = 16'h0000;
	mel_filter_coefs[19][96] = 16'h0000;
	mel_filter_coefs[19][97] = 16'h0000;
	mel_filter_coefs[19][98] = 16'h0000;
	mel_filter_coefs[19][99] = 16'h0000;
	mel_filter_coefs[19][100] = 16'h0000;
	mel_filter_coefs[19][101] = 16'h0000;
	mel_filter_coefs[19][102] = 16'h0000;
	mel_filter_coefs[19][103] = 16'h0000;
	mel_filter_coefs[19][104] = 16'h0000;
	mel_filter_coefs[19][105] = 16'h0000;
	mel_filter_coefs[19][106] = 16'h0000;
	mel_filter_coefs[19][107] = 16'h0000;
	mel_filter_coefs[19][108] = 16'h0000;
	mel_filter_coefs[19][109] = 16'h0000;
	mel_filter_coefs[19][110] = 16'h0000;
	mel_filter_coefs[19][111] = 16'h0000;
	mel_filter_coefs[19][112] = 16'h0000;
	mel_filter_coefs[19][113] = 16'h0000;
	mel_filter_coefs[19][114] = 16'h0000;
	mel_filter_coefs[19][115] = 16'h0000;
	mel_filter_coefs[19][116] = 16'h0000;
	mel_filter_coefs[19][117] = 16'h0000;
	mel_filter_coefs[19][118] = 16'h0000;
	mel_filter_coefs[19][119] = 16'h0000;
	mel_filter_coefs[19][120] = 16'h0000;
	mel_filter_coefs[19][121] = 16'h0000;
	mel_filter_coefs[19][122] = 16'h0000;
	mel_filter_coefs[19][123] = 16'h0000;
	mel_filter_coefs[19][124] = 16'h0000;
	mel_filter_coefs[19][125] = 16'h0000;
	mel_filter_coefs[19][126] = 16'h0000;
	mel_filter_coefs[19][127] = 16'h0000;
	mel_filter_coefs[19][128] = 16'h0000;
	mel_filter_coefs[19][129] = 16'h0000;
	mel_filter_coefs[19][130] = 16'h0000;
	mel_filter_coefs[19][131] = 16'h0000;
	mel_filter_coefs[19][132] = 16'h0000;
	mel_filter_coefs[19][133] = 16'h0000;
	mel_filter_coefs[19][134] = 16'h0000;
	mel_filter_coefs[19][135] = 16'h0000;
	mel_filter_coefs[19][136] = 16'h0000;
	mel_filter_coefs[19][137] = 16'h0000;
	mel_filter_coefs[19][138] = 16'h0000;
	mel_filter_coefs[19][139] = 16'h0000;
	mel_filter_coefs[19][140] = 16'h0000;
	mel_filter_coefs[19][141] = 16'h0000;
	mel_filter_coefs[19][142] = 16'h0000;
	mel_filter_coefs[19][143] = 16'h0000;
	mel_filter_coefs[19][144] = 16'h0000;
	mel_filter_coefs[19][145] = 16'h0000;
	mel_filter_coefs[19][146] = 16'h0000;
	mel_filter_coefs[19][147] = 16'h0000;
	mel_filter_coefs[19][148] = 16'h0000;
	mel_filter_coefs[19][149] = 16'h0000;
	mel_filter_coefs[19][150] = 16'h0000;
	mel_filter_coefs[19][151] = 16'h0000;
	mel_filter_coefs[19][152] = 16'h0000;
	mel_filter_coefs[19][153] = 16'h0000;
	mel_filter_coefs[19][154] = 16'h0000;
	mel_filter_coefs[19][155] = 16'h0000;
	mel_filter_coefs[19][156] = 16'h0000;
	mel_filter_coefs[19][157] = 16'h0000;
	mel_filter_coefs[19][158] = 16'h0000;
	mel_filter_coefs[19][159] = 16'h0000;
	mel_filter_coefs[19][160] = 16'h0000;
	mel_filter_coefs[19][161] = 16'h0000;
	mel_filter_coefs[19][162] = 16'h0000;
	mel_filter_coefs[19][163] = 16'h0000;
	mel_filter_coefs[19][164] = 16'h0000;
	mel_filter_coefs[19][165] = 16'h0000;
	mel_filter_coefs[19][166] = 16'h0000;
	mel_filter_coefs[19][167] = 16'h0000;
	mel_filter_coefs[19][168] = 16'h0000;
	mel_filter_coefs[19][169] = 16'h0000;
	mel_filter_coefs[19][170] = 16'h0000;
	mel_filter_coefs[19][171] = 16'h0000;
	mel_filter_coefs[19][172] = 16'h0000;
	mel_filter_coefs[19][173] = 16'h0000;
	mel_filter_coefs[19][174] = 16'h0000;
	mel_filter_coefs[19][175] = 16'h0000;
	mel_filter_coefs[19][176] = 16'h0000;
	mel_filter_coefs[19][177] = 16'h0000;
	mel_filter_coefs[19][178] = 16'h0000;
	mel_filter_coefs[19][179] = 16'h0000;
	mel_filter_coefs[19][180] = 16'h0000;
	mel_filter_coefs[19][181] = 16'h0000;
	mel_filter_coefs[19][182] = 16'h0000;
	mel_filter_coefs[19][183] = 16'h0000;
	mel_filter_coefs[19][184] = 16'h0000;
	mel_filter_coefs[19][185] = 16'h0000;
	mel_filter_coefs[19][186] = 16'h0000;
	mel_filter_coefs[19][187] = 16'h0000;
	mel_filter_coefs[19][188] = 16'h0000;
	mel_filter_coefs[19][189] = 16'h0000;
	mel_filter_coefs[19][190] = 16'h0000;
	mel_filter_coefs[19][191] = 16'h0000;
	mel_filter_coefs[19][192] = 16'h0000;
	mel_filter_coefs[19][193] = 16'h0000;
	mel_filter_coefs[19][194] = 16'h0000;
	mel_filter_coefs[19][195] = 16'h0000;
	mel_filter_coefs[19][196] = 16'h0000;
	mel_filter_coefs[19][197] = 16'h0000;
	mel_filter_coefs[19][198] = 16'h0000;
	mel_filter_coefs[19][199] = 16'h0000;
	mel_filter_coefs[19][200] = 16'h0000;
	mel_filter_coefs[19][201] = 16'h0000;
	mel_filter_coefs[19][202] = 16'h0000;
	mel_filter_coefs[19][203] = 16'h0000;
	mel_filter_coefs[19][204] = 16'h0000;
	mel_filter_coefs[19][205] = 16'h0000;
	mel_filter_coefs[19][206] = 16'h0000;
	mel_filter_coefs[19][207] = 16'h0000;
	mel_filter_coefs[19][208] = 16'h0000;
	mel_filter_coefs[19][209] = 16'h0000;
	mel_filter_coefs[19][210] = 16'h0000;
	mel_filter_coefs[19][211] = 16'h0000;
	mel_filter_coefs[19][212] = 16'h0000;
	mel_filter_coefs[19][213] = 16'h0000;
	mel_filter_coefs[19][214] = 16'h0000;
	mel_filter_coefs[19][215] = 16'h0000;
	mel_filter_coefs[19][216] = 16'h0000;
	mel_filter_coefs[19][217] = 16'h0000;
	mel_filter_coefs[19][218] = 16'h0000;
	mel_filter_coefs[19][219] = 16'h0000;
	mel_filter_coefs[19][220] = 16'h0000;
	mel_filter_coefs[19][221] = 16'h0000;
	mel_filter_coefs[19][222] = 16'h0000;
	mel_filter_coefs[19][223] = 16'h0000;
	mel_filter_coefs[19][224] = 16'h0000;
	mel_filter_coefs[19][225] = 16'h0000;
	mel_filter_coefs[19][226] = 16'h0000;
	mel_filter_coefs[19][227] = 16'h0000;
	mel_filter_coefs[19][228] = 16'h0000;
	mel_filter_coefs[19][229] = 16'h0000;
	mel_filter_coefs[19][230] = 16'h0000;
	mel_filter_coefs[19][231] = 16'h0000;
	mel_filter_coefs[19][232] = 16'h0000;
	mel_filter_coefs[19][233] = 16'h0000;
	mel_filter_coefs[19][234] = 16'h0000;
	mel_filter_coefs[19][235] = 16'h0000;
	mel_filter_coefs[19][236] = 16'h0000;
	mel_filter_coefs[19][237] = 16'h0000;
	mel_filter_coefs[19][238] = 16'h0000;
	mel_filter_coefs[19][239] = 16'h0000;
	mel_filter_coefs[19][240] = 16'h0000;
	mel_filter_coefs[19][241] = 16'h0000;
	mel_filter_coefs[19][242] = 16'h0000;
	mel_filter_coefs[19][243] = 16'h0000;
	mel_filter_coefs[19][244] = 16'h0000;
	mel_filter_coefs[19][245] = 16'h0000;
	mel_filter_coefs[19][246] = 16'h0000;
	mel_filter_coefs[19][247] = 16'h0000;
	mel_filter_coefs[19][248] = 16'h0000;
	mel_filter_coefs[19][249] = 16'h0000;
	mel_filter_coefs[19][250] = 16'h0000;
	mel_filter_coefs[19][251] = 16'h0000;
	mel_filter_coefs[19][252] = 16'h0000;
	mel_filter_coefs[19][253] = 16'h0000;
	mel_filter_coefs[19][254] = 16'h0000;
	mel_filter_coefs[19][255] = 16'h0000;
	mel_filter_coefs[20][0] = 16'h0000;
	mel_filter_coefs[20][1] = 16'h0000;
	mel_filter_coefs[20][2] = 16'h0000;
	mel_filter_coefs[20][3] = 16'h0000;
	mel_filter_coefs[20][4] = 16'h0000;
	mel_filter_coefs[20][5] = 16'h0000;
	mel_filter_coefs[20][6] = 16'h0000;
	mel_filter_coefs[20][7] = 16'h0000;
	mel_filter_coefs[20][8] = 16'h0000;
	mel_filter_coefs[20][9] = 16'h0000;
	mel_filter_coefs[20][10] = 16'h0000;
	mel_filter_coefs[20][11] = 16'h0000;
	mel_filter_coefs[20][12] = 16'h0000;
	mel_filter_coefs[20][13] = 16'h0000;
	mel_filter_coefs[20][14] = 16'h0000;
	mel_filter_coefs[20][15] = 16'h0000;
	mel_filter_coefs[20][16] = 16'h0000;
	mel_filter_coefs[20][17] = 16'h0000;
	mel_filter_coefs[20][18] = 16'h0000;
	mel_filter_coefs[20][19] = 16'h0000;
	mel_filter_coefs[20][20] = 16'h0000;
	mel_filter_coefs[20][21] = 16'h0000;
	mel_filter_coefs[20][22] = 16'h0000;
	mel_filter_coefs[20][23] = 16'h0000;
	mel_filter_coefs[20][24] = 16'h0000;
	mel_filter_coefs[20][25] = 16'h0000;
	mel_filter_coefs[20][26] = 16'h0000;
	mel_filter_coefs[20][27] = 16'h0000;
	mel_filter_coefs[20][28] = 16'h0000;
	mel_filter_coefs[20][29] = 16'h0000;
	mel_filter_coefs[20][30] = 16'h0000;
	mel_filter_coefs[20][31] = 16'h0000;
	mel_filter_coefs[20][32] = 16'h0000;
	mel_filter_coefs[20][33] = 16'h0000;
	mel_filter_coefs[20][34] = 16'h0000;
	mel_filter_coefs[20][35] = 16'h0000;
	mel_filter_coefs[20][36] = 16'h0000;
	mel_filter_coefs[20][37] = 16'h0000;
	mel_filter_coefs[20][38] = 16'h0000;
	mel_filter_coefs[20][39] = 16'h0000;
	mel_filter_coefs[20][40] = 16'h0000;
	mel_filter_coefs[20][41] = 16'h0000;
	mel_filter_coefs[20][42] = 16'h0000;
	mel_filter_coefs[20][43] = 16'h0000;
	mel_filter_coefs[20][44] = 16'h0000;
	mel_filter_coefs[20][45] = 16'h0000;
	mel_filter_coefs[20][46] = 16'h0000;
	mel_filter_coefs[20][47] = 16'h0000;
	mel_filter_coefs[20][48] = 16'h0000;
	mel_filter_coefs[20][49] = 16'h0000;
	mel_filter_coefs[20][50] = 16'h0000;
	mel_filter_coefs[20][51] = 16'h0000;
	mel_filter_coefs[20][52] = 16'h0000;
	mel_filter_coefs[20][53] = 16'h0000;
	mel_filter_coefs[20][54] = 16'h00DA;
	mel_filter_coefs[20][55] = 16'h1B53;
	mel_filter_coefs[20][56] = 16'h35CB;
	mel_filter_coefs[20][57] = 16'h5044;
	mel_filter_coefs[20][58] = 16'h6ABC;
	mel_filter_coefs[20][59] = 16'h7B1B;
	mel_filter_coefs[20][60] = 16'h6236;
	mel_filter_coefs[20][61] = 16'h4951;
	mel_filter_coefs[20][62] = 16'h306D;
	mel_filter_coefs[20][63] = 16'h1788;
	mel_filter_coefs[20][64] = 16'h0000;
	mel_filter_coefs[20][65] = 16'h0000;
	mel_filter_coefs[20][66] = 16'h0000;
	mel_filter_coefs[20][67] = 16'h0000;
	mel_filter_coefs[20][68] = 16'h0000;
	mel_filter_coefs[20][69] = 16'h0000;
	mel_filter_coefs[20][70] = 16'h0000;
	mel_filter_coefs[20][71] = 16'h0000;
	mel_filter_coefs[20][72] = 16'h0000;
	mel_filter_coefs[20][73] = 16'h0000;
	mel_filter_coefs[20][74] = 16'h0000;
	mel_filter_coefs[20][75] = 16'h0000;
	mel_filter_coefs[20][76] = 16'h0000;
	mel_filter_coefs[20][77] = 16'h0000;
	mel_filter_coefs[20][78] = 16'h0000;
	mel_filter_coefs[20][79] = 16'h0000;
	mel_filter_coefs[20][80] = 16'h0000;
	mel_filter_coefs[20][81] = 16'h0000;
	mel_filter_coefs[20][82] = 16'h0000;
	mel_filter_coefs[20][83] = 16'h0000;
	mel_filter_coefs[20][84] = 16'h0000;
	mel_filter_coefs[20][85] = 16'h0000;
	mel_filter_coefs[20][86] = 16'h0000;
	mel_filter_coefs[20][87] = 16'h0000;
	mel_filter_coefs[20][88] = 16'h0000;
	mel_filter_coefs[20][89] = 16'h0000;
	mel_filter_coefs[20][90] = 16'h0000;
	mel_filter_coefs[20][91] = 16'h0000;
	mel_filter_coefs[20][92] = 16'h0000;
	mel_filter_coefs[20][93] = 16'h0000;
	mel_filter_coefs[20][94] = 16'h0000;
	mel_filter_coefs[20][95] = 16'h0000;
	mel_filter_coefs[20][96] = 16'h0000;
	mel_filter_coefs[20][97] = 16'h0000;
	mel_filter_coefs[20][98] = 16'h0000;
	mel_filter_coefs[20][99] = 16'h0000;
	mel_filter_coefs[20][100] = 16'h0000;
	mel_filter_coefs[20][101] = 16'h0000;
	mel_filter_coefs[20][102] = 16'h0000;
	mel_filter_coefs[20][103] = 16'h0000;
	mel_filter_coefs[20][104] = 16'h0000;
	mel_filter_coefs[20][105] = 16'h0000;
	mel_filter_coefs[20][106] = 16'h0000;
	mel_filter_coefs[20][107] = 16'h0000;
	mel_filter_coefs[20][108] = 16'h0000;
	mel_filter_coefs[20][109] = 16'h0000;
	mel_filter_coefs[20][110] = 16'h0000;
	mel_filter_coefs[20][111] = 16'h0000;
	mel_filter_coefs[20][112] = 16'h0000;
	mel_filter_coefs[20][113] = 16'h0000;
	mel_filter_coefs[20][114] = 16'h0000;
	mel_filter_coefs[20][115] = 16'h0000;
	mel_filter_coefs[20][116] = 16'h0000;
	mel_filter_coefs[20][117] = 16'h0000;
	mel_filter_coefs[20][118] = 16'h0000;
	mel_filter_coefs[20][119] = 16'h0000;
	mel_filter_coefs[20][120] = 16'h0000;
	mel_filter_coefs[20][121] = 16'h0000;
	mel_filter_coefs[20][122] = 16'h0000;
	mel_filter_coefs[20][123] = 16'h0000;
	mel_filter_coefs[20][124] = 16'h0000;
	mel_filter_coefs[20][125] = 16'h0000;
	mel_filter_coefs[20][126] = 16'h0000;
	mel_filter_coefs[20][127] = 16'h0000;
	mel_filter_coefs[20][128] = 16'h0000;
	mel_filter_coefs[20][129] = 16'h0000;
	mel_filter_coefs[20][130] = 16'h0000;
	mel_filter_coefs[20][131] = 16'h0000;
	mel_filter_coefs[20][132] = 16'h0000;
	mel_filter_coefs[20][133] = 16'h0000;
	mel_filter_coefs[20][134] = 16'h0000;
	mel_filter_coefs[20][135] = 16'h0000;
	mel_filter_coefs[20][136] = 16'h0000;
	mel_filter_coefs[20][137] = 16'h0000;
	mel_filter_coefs[20][138] = 16'h0000;
	mel_filter_coefs[20][139] = 16'h0000;
	mel_filter_coefs[20][140] = 16'h0000;
	mel_filter_coefs[20][141] = 16'h0000;
	mel_filter_coefs[20][142] = 16'h0000;
	mel_filter_coefs[20][143] = 16'h0000;
	mel_filter_coefs[20][144] = 16'h0000;
	mel_filter_coefs[20][145] = 16'h0000;
	mel_filter_coefs[20][146] = 16'h0000;
	mel_filter_coefs[20][147] = 16'h0000;
	mel_filter_coefs[20][148] = 16'h0000;
	mel_filter_coefs[20][149] = 16'h0000;
	mel_filter_coefs[20][150] = 16'h0000;
	mel_filter_coefs[20][151] = 16'h0000;
	mel_filter_coefs[20][152] = 16'h0000;
	mel_filter_coefs[20][153] = 16'h0000;
	mel_filter_coefs[20][154] = 16'h0000;
	mel_filter_coefs[20][155] = 16'h0000;
	mel_filter_coefs[20][156] = 16'h0000;
	mel_filter_coefs[20][157] = 16'h0000;
	mel_filter_coefs[20][158] = 16'h0000;
	mel_filter_coefs[20][159] = 16'h0000;
	mel_filter_coefs[20][160] = 16'h0000;
	mel_filter_coefs[20][161] = 16'h0000;
	mel_filter_coefs[20][162] = 16'h0000;
	mel_filter_coefs[20][163] = 16'h0000;
	mel_filter_coefs[20][164] = 16'h0000;
	mel_filter_coefs[20][165] = 16'h0000;
	mel_filter_coefs[20][166] = 16'h0000;
	mel_filter_coefs[20][167] = 16'h0000;
	mel_filter_coefs[20][168] = 16'h0000;
	mel_filter_coefs[20][169] = 16'h0000;
	mel_filter_coefs[20][170] = 16'h0000;
	mel_filter_coefs[20][171] = 16'h0000;
	mel_filter_coefs[20][172] = 16'h0000;
	mel_filter_coefs[20][173] = 16'h0000;
	mel_filter_coefs[20][174] = 16'h0000;
	mel_filter_coefs[20][175] = 16'h0000;
	mel_filter_coefs[20][176] = 16'h0000;
	mel_filter_coefs[20][177] = 16'h0000;
	mel_filter_coefs[20][178] = 16'h0000;
	mel_filter_coefs[20][179] = 16'h0000;
	mel_filter_coefs[20][180] = 16'h0000;
	mel_filter_coefs[20][181] = 16'h0000;
	mel_filter_coefs[20][182] = 16'h0000;
	mel_filter_coefs[20][183] = 16'h0000;
	mel_filter_coefs[20][184] = 16'h0000;
	mel_filter_coefs[20][185] = 16'h0000;
	mel_filter_coefs[20][186] = 16'h0000;
	mel_filter_coefs[20][187] = 16'h0000;
	mel_filter_coefs[20][188] = 16'h0000;
	mel_filter_coefs[20][189] = 16'h0000;
	mel_filter_coefs[20][190] = 16'h0000;
	mel_filter_coefs[20][191] = 16'h0000;
	mel_filter_coefs[20][192] = 16'h0000;
	mel_filter_coefs[20][193] = 16'h0000;
	mel_filter_coefs[20][194] = 16'h0000;
	mel_filter_coefs[20][195] = 16'h0000;
	mel_filter_coefs[20][196] = 16'h0000;
	mel_filter_coefs[20][197] = 16'h0000;
	mel_filter_coefs[20][198] = 16'h0000;
	mel_filter_coefs[20][199] = 16'h0000;
	mel_filter_coefs[20][200] = 16'h0000;
	mel_filter_coefs[20][201] = 16'h0000;
	mel_filter_coefs[20][202] = 16'h0000;
	mel_filter_coefs[20][203] = 16'h0000;
	mel_filter_coefs[20][204] = 16'h0000;
	mel_filter_coefs[20][205] = 16'h0000;
	mel_filter_coefs[20][206] = 16'h0000;
	mel_filter_coefs[20][207] = 16'h0000;
	mel_filter_coefs[20][208] = 16'h0000;
	mel_filter_coefs[20][209] = 16'h0000;
	mel_filter_coefs[20][210] = 16'h0000;
	mel_filter_coefs[20][211] = 16'h0000;
	mel_filter_coefs[20][212] = 16'h0000;
	mel_filter_coefs[20][213] = 16'h0000;
	mel_filter_coefs[20][214] = 16'h0000;
	mel_filter_coefs[20][215] = 16'h0000;
	mel_filter_coefs[20][216] = 16'h0000;
	mel_filter_coefs[20][217] = 16'h0000;
	mel_filter_coefs[20][218] = 16'h0000;
	mel_filter_coefs[20][219] = 16'h0000;
	mel_filter_coefs[20][220] = 16'h0000;
	mel_filter_coefs[20][221] = 16'h0000;
	mel_filter_coefs[20][222] = 16'h0000;
	mel_filter_coefs[20][223] = 16'h0000;
	mel_filter_coefs[20][224] = 16'h0000;
	mel_filter_coefs[20][225] = 16'h0000;
	mel_filter_coefs[20][226] = 16'h0000;
	mel_filter_coefs[20][227] = 16'h0000;
	mel_filter_coefs[20][228] = 16'h0000;
	mel_filter_coefs[20][229] = 16'h0000;
	mel_filter_coefs[20][230] = 16'h0000;
	mel_filter_coefs[20][231] = 16'h0000;
	mel_filter_coefs[20][232] = 16'h0000;
	mel_filter_coefs[20][233] = 16'h0000;
	mel_filter_coefs[20][234] = 16'h0000;
	mel_filter_coefs[20][235] = 16'h0000;
	mel_filter_coefs[20][236] = 16'h0000;
	mel_filter_coefs[20][237] = 16'h0000;
	mel_filter_coefs[20][238] = 16'h0000;
	mel_filter_coefs[20][239] = 16'h0000;
	mel_filter_coefs[20][240] = 16'h0000;
	mel_filter_coefs[20][241] = 16'h0000;
	mel_filter_coefs[20][242] = 16'h0000;
	mel_filter_coefs[20][243] = 16'h0000;
	mel_filter_coefs[20][244] = 16'h0000;
	mel_filter_coefs[20][245] = 16'h0000;
	mel_filter_coefs[20][246] = 16'h0000;
	mel_filter_coefs[20][247] = 16'h0000;
	mel_filter_coefs[20][248] = 16'h0000;
	mel_filter_coefs[20][249] = 16'h0000;
	mel_filter_coefs[20][250] = 16'h0000;
	mel_filter_coefs[20][251] = 16'h0000;
	mel_filter_coefs[20][252] = 16'h0000;
	mel_filter_coefs[20][253] = 16'h0000;
	mel_filter_coefs[20][254] = 16'h0000;
	mel_filter_coefs[20][255] = 16'h0000;
	mel_filter_coefs[21][0] = 16'h0000;
	mel_filter_coefs[21][1] = 16'h0000;
	mel_filter_coefs[21][2] = 16'h0000;
	mel_filter_coefs[21][3] = 16'h0000;
	mel_filter_coefs[21][4] = 16'h0000;
	mel_filter_coefs[21][5] = 16'h0000;
	mel_filter_coefs[21][6] = 16'h0000;
	mel_filter_coefs[21][7] = 16'h0000;
	mel_filter_coefs[21][8] = 16'h0000;
	mel_filter_coefs[21][9] = 16'h0000;
	mel_filter_coefs[21][10] = 16'h0000;
	mel_filter_coefs[21][11] = 16'h0000;
	mel_filter_coefs[21][12] = 16'h0000;
	mel_filter_coefs[21][13] = 16'h0000;
	mel_filter_coefs[21][14] = 16'h0000;
	mel_filter_coefs[21][15] = 16'h0000;
	mel_filter_coefs[21][16] = 16'h0000;
	mel_filter_coefs[21][17] = 16'h0000;
	mel_filter_coefs[21][18] = 16'h0000;
	mel_filter_coefs[21][19] = 16'h0000;
	mel_filter_coefs[21][20] = 16'h0000;
	mel_filter_coefs[21][21] = 16'h0000;
	mel_filter_coefs[21][22] = 16'h0000;
	mel_filter_coefs[21][23] = 16'h0000;
	mel_filter_coefs[21][24] = 16'h0000;
	mel_filter_coefs[21][25] = 16'h0000;
	mel_filter_coefs[21][26] = 16'h0000;
	mel_filter_coefs[21][27] = 16'h0000;
	mel_filter_coefs[21][28] = 16'h0000;
	mel_filter_coefs[21][29] = 16'h0000;
	mel_filter_coefs[21][30] = 16'h0000;
	mel_filter_coefs[21][31] = 16'h0000;
	mel_filter_coefs[21][32] = 16'h0000;
	mel_filter_coefs[21][33] = 16'h0000;
	mel_filter_coefs[21][34] = 16'h0000;
	mel_filter_coefs[21][35] = 16'h0000;
	mel_filter_coefs[21][36] = 16'h0000;
	mel_filter_coefs[21][37] = 16'h0000;
	mel_filter_coefs[21][38] = 16'h0000;
	mel_filter_coefs[21][39] = 16'h0000;
	mel_filter_coefs[21][40] = 16'h0000;
	mel_filter_coefs[21][41] = 16'h0000;
	mel_filter_coefs[21][42] = 16'h0000;
	mel_filter_coefs[21][43] = 16'h0000;
	mel_filter_coefs[21][44] = 16'h0000;
	mel_filter_coefs[21][45] = 16'h0000;
	mel_filter_coefs[21][46] = 16'h0000;
	mel_filter_coefs[21][47] = 16'h0000;
	mel_filter_coefs[21][48] = 16'h0000;
	mel_filter_coefs[21][49] = 16'h0000;
	mel_filter_coefs[21][50] = 16'h0000;
	mel_filter_coefs[21][51] = 16'h0000;
	mel_filter_coefs[21][52] = 16'h0000;
	mel_filter_coefs[21][53] = 16'h0000;
	mel_filter_coefs[21][54] = 16'h0000;
	mel_filter_coefs[21][55] = 16'h0000;
	mel_filter_coefs[21][56] = 16'h0000;
	mel_filter_coefs[21][57] = 16'h0000;
	mel_filter_coefs[21][58] = 16'h0000;
	mel_filter_coefs[21][59] = 16'h04E5;
	mel_filter_coefs[21][60] = 16'h1DCA;
	mel_filter_coefs[21][61] = 16'h36AF;
	mel_filter_coefs[21][62] = 16'h4F93;
	mel_filter_coefs[21][63] = 16'h6878;
	mel_filter_coefs[21][64] = 16'h7EB9;
	mel_filter_coefs[21][65] = 16'h6750;
	mel_filter_coefs[21][66] = 16'h4FE7;
	mel_filter_coefs[21][67] = 16'h387F;
	mel_filter_coefs[21][68] = 16'h2116;
	mel_filter_coefs[21][69] = 16'h09AD;
	mel_filter_coefs[21][70] = 16'h0000;
	mel_filter_coefs[21][71] = 16'h0000;
	mel_filter_coefs[21][72] = 16'h0000;
	mel_filter_coefs[21][73] = 16'h0000;
	mel_filter_coefs[21][74] = 16'h0000;
	mel_filter_coefs[21][75] = 16'h0000;
	mel_filter_coefs[21][76] = 16'h0000;
	mel_filter_coefs[21][77] = 16'h0000;
	mel_filter_coefs[21][78] = 16'h0000;
	mel_filter_coefs[21][79] = 16'h0000;
	mel_filter_coefs[21][80] = 16'h0000;
	mel_filter_coefs[21][81] = 16'h0000;
	mel_filter_coefs[21][82] = 16'h0000;
	mel_filter_coefs[21][83] = 16'h0000;
	mel_filter_coefs[21][84] = 16'h0000;
	mel_filter_coefs[21][85] = 16'h0000;
	mel_filter_coefs[21][86] = 16'h0000;
	mel_filter_coefs[21][87] = 16'h0000;
	mel_filter_coefs[21][88] = 16'h0000;
	mel_filter_coefs[21][89] = 16'h0000;
	mel_filter_coefs[21][90] = 16'h0000;
	mel_filter_coefs[21][91] = 16'h0000;
	mel_filter_coefs[21][92] = 16'h0000;
	mel_filter_coefs[21][93] = 16'h0000;
	mel_filter_coefs[21][94] = 16'h0000;
	mel_filter_coefs[21][95] = 16'h0000;
	mel_filter_coefs[21][96] = 16'h0000;
	mel_filter_coefs[21][97] = 16'h0000;
	mel_filter_coefs[21][98] = 16'h0000;
	mel_filter_coefs[21][99] = 16'h0000;
	mel_filter_coefs[21][100] = 16'h0000;
	mel_filter_coefs[21][101] = 16'h0000;
	mel_filter_coefs[21][102] = 16'h0000;
	mel_filter_coefs[21][103] = 16'h0000;
	mel_filter_coefs[21][104] = 16'h0000;
	mel_filter_coefs[21][105] = 16'h0000;
	mel_filter_coefs[21][106] = 16'h0000;
	mel_filter_coefs[21][107] = 16'h0000;
	mel_filter_coefs[21][108] = 16'h0000;
	mel_filter_coefs[21][109] = 16'h0000;
	mel_filter_coefs[21][110] = 16'h0000;
	mel_filter_coefs[21][111] = 16'h0000;
	mel_filter_coefs[21][112] = 16'h0000;
	mel_filter_coefs[21][113] = 16'h0000;
	mel_filter_coefs[21][114] = 16'h0000;
	mel_filter_coefs[21][115] = 16'h0000;
	mel_filter_coefs[21][116] = 16'h0000;
	mel_filter_coefs[21][117] = 16'h0000;
	mel_filter_coefs[21][118] = 16'h0000;
	mel_filter_coefs[21][119] = 16'h0000;
	mel_filter_coefs[21][120] = 16'h0000;
	mel_filter_coefs[21][121] = 16'h0000;
	mel_filter_coefs[21][122] = 16'h0000;
	mel_filter_coefs[21][123] = 16'h0000;
	mel_filter_coefs[21][124] = 16'h0000;
	mel_filter_coefs[21][125] = 16'h0000;
	mel_filter_coefs[21][126] = 16'h0000;
	mel_filter_coefs[21][127] = 16'h0000;
	mel_filter_coefs[21][128] = 16'h0000;
	mel_filter_coefs[21][129] = 16'h0000;
	mel_filter_coefs[21][130] = 16'h0000;
	mel_filter_coefs[21][131] = 16'h0000;
	mel_filter_coefs[21][132] = 16'h0000;
	mel_filter_coefs[21][133] = 16'h0000;
	mel_filter_coefs[21][134] = 16'h0000;
	mel_filter_coefs[21][135] = 16'h0000;
	mel_filter_coefs[21][136] = 16'h0000;
	mel_filter_coefs[21][137] = 16'h0000;
	mel_filter_coefs[21][138] = 16'h0000;
	mel_filter_coefs[21][139] = 16'h0000;
	mel_filter_coefs[21][140] = 16'h0000;
	mel_filter_coefs[21][141] = 16'h0000;
	mel_filter_coefs[21][142] = 16'h0000;
	mel_filter_coefs[21][143] = 16'h0000;
	mel_filter_coefs[21][144] = 16'h0000;
	mel_filter_coefs[21][145] = 16'h0000;
	mel_filter_coefs[21][146] = 16'h0000;
	mel_filter_coefs[21][147] = 16'h0000;
	mel_filter_coefs[21][148] = 16'h0000;
	mel_filter_coefs[21][149] = 16'h0000;
	mel_filter_coefs[21][150] = 16'h0000;
	mel_filter_coefs[21][151] = 16'h0000;
	mel_filter_coefs[21][152] = 16'h0000;
	mel_filter_coefs[21][153] = 16'h0000;
	mel_filter_coefs[21][154] = 16'h0000;
	mel_filter_coefs[21][155] = 16'h0000;
	mel_filter_coefs[21][156] = 16'h0000;
	mel_filter_coefs[21][157] = 16'h0000;
	mel_filter_coefs[21][158] = 16'h0000;
	mel_filter_coefs[21][159] = 16'h0000;
	mel_filter_coefs[21][160] = 16'h0000;
	mel_filter_coefs[21][161] = 16'h0000;
	mel_filter_coefs[21][162] = 16'h0000;
	mel_filter_coefs[21][163] = 16'h0000;
	mel_filter_coefs[21][164] = 16'h0000;
	mel_filter_coefs[21][165] = 16'h0000;
	mel_filter_coefs[21][166] = 16'h0000;
	mel_filter_coefs[21][167] = 16'h0000;
	mel_filter_coefs[21][168] = 16'h0000;
	mel_filter_coefs[21][169] = 16'h0000;
	mel_filter_coefs[21][170] = 16'h0000;
	mel_filter_coefs[21][171] = 16'h0000;
	mel_filter_coefs[21][172] = 16'h0000;
	mel_filter_coefs[21][173] = 16'h0000;
	mel_filter_coefs[21][174] = 16'h0000;
	mel_filter_coefs[21][175] = 16'h0000;
	mel_filter_coefs[21][176] = 16'h0000;
	mel_filter_coefs[21][177] = 16'h0000;
	mel_filter_coefs[21][178] = 16'h0000;
	mel_filter_coefs[21][179] = 16'h0000;
	mel_filter_coefs[21][180] = 16'h0000;
	mel_filter_coefs[21][181] = 16'h0000;
	mel_filter_coefs[21][182] = 16'h0000;
	mel_filter_coefs[21][183] = 16'h0000;
	mel_filter_coefs[21][184] = 16'h0000;
	mel_filter_coefs[21][185] = 16'h0000;
	mel_filter_coefs[21][186] = 16'h0000;
	mel_filter_coefs[21][187] = 16'h0000;
	mel_filter_coefs[21][188] = 16'h0000;
	mel_filter_coefs[21][189] = 16'h0000;
	mel_filter_coefs[21][190] = 16'h0000;
	mel_filter_coefs[21][191] = 16'h0000;
	mel_filter_coefs[21][192] = 16'h0000;
	mel_filter_coefs[21][193] = 16'h0000;
	mel_filter_coefs[21][194] = 16'h0000;
	mel_filter_coefs[21][195] = 16'h0000;
	mel_filter_coefs[21][196] = 16'h0000;
	mel_filter_coefs[21][197] = 16'h0000;
	mel_filter_coefs[21][198] = 16'h0000;
	mel_filter_coefs[21][199] = 16'h0000;
	mel_filter_coefs[21][200] = 16'h0000;
	mel_filter_coefs[21][201] = 16'h0000;
	mel_filter_coefs[21][202] = 16'h0000;
	mel_filter_coefs[21][203] = 16'h0000;
	mel_filter_coefs[21][204] = 16'h0000;
	mel_filter_coefs[21][205] = 16'h0000;
	mel_filter_coefs[21][206] = 16'h0000;
	mel_filter_coefs[21][207] = 16'h0000;
	mel_filter_coefs[21][208] = 16'h0000;
	mel_filter_coefs[21][209] = 16'h0000;
	mel_filter_coefs[21][210] = 16'h0000;
	mel_filter_coefs[21][211] = 16'h0000;
	mel_filter_coefs[21][212] = 16'h0000;
	mel_filter_coefs[21][213] = 16'h0000;
	mel_filter_coefs[21][214] = 16'h0000;
	mel_filter_coefs[21][215] = 16'h0000;
	mel_filter_coefs[21][216] = 16'h0000;
	mel_filter_coefs[21][217] = 16'h0000;
	mel_filter_coefs[21][218] = 16'h0000;
	mel_filter_coefs[21][219] = 16'h0000;
	mel_filter_coefs[21][220] = 16'h0000;
	mel_filter_coefs[21][221] = 16'h0000;
	mel_filter_coefs[21][222] = 16'h0000;
	mel_filter_coefs[21][223] = 16'h0000;
	mel_filter_coefs[21][224] = 16'h0000;
	mel_filter_coefs[21][225] = 16'h0000;
	mel_filter_coefs[21][226] = 16'h0000;
	mel_filter_coefs[21][227] = 16'h0000;
	mel_filter_coefs[21][228] = 16'h0000;
	mel_filter_coefs[21][229] = 16'h0000;
	mel_filter_coefs[21][230] = 16'h0000;
	mel_filter_coefs[21][231] = 16'h0000;
	mel_filter_coefs[21][232] = 16'h0000;
	mel_filter_coefs[21][233] = 16'h0000;
	mel_filter_coefs[21][234] = 16'h0000;
	mel_filter_coefs[21][235] = 16'h0000;
	mel_filter_coefs[21][236] = 16'h0000;
	mel_filter_coefs[21][237] = 16'h0000;
	mel_filter_coefs[21][238] = 16'h0000;
	mel_filter_coefs[21][239] = 16'h0000;
	mel_filter_coefs[21][240] = 16'h0000;
	mel_filter_coefs[21][241] = 16'h0000;
	mel_filter_coefs[21][242] = 16'h0000;
	mel_filter_coefs[21][243] = 16'h0000;
	mel_filter_coefs[21][244] = 16'h0000;
	mel_filter_coefs[21][245] = 16'h0000;
	mel_filter_coefs[21][246] = 16'h0000;
	mel_filter_coefs[21][247] = 16'h0000;
	mel_filter_coefs[21][248] = 16'h0000;
	mel_filter_coefs[21][249] = 16'h0000;
	mel_filter_coefs[21][250] = 16'h0000;
	mel_filter_coefs[21][251] = 16'h0000;
	mel_filter_coefs[21][252] = 16'h0000;
	mel_filter_coefs[21][253] = 16'h0000;
	mel_filter_coefs[21][254] = 16'h0000;
	mel_filter_coefs[21][255] = 16'h0000;
	mel_filter_coefs[22][0] = 16'h0000;
	mel_filter_coefs[22][1] = 16'h0000;
	mel_filter_coefs[22][2] = 16'h0000;
	mel_filter_coefs[22][3] = 16'h0000;
	mel_filter_coefs[22][4] = 16'h0000;
	mel_filter_coefs[22][5] = 16'h0000;
	mel_filter_coefs[22][6] = 16'h0000;
	mel_filter_coefs[22][7] = 16'h0000;
	mel_filter_coefs[22][8] = 16'h0000;
	mel_filter_coefs[22][9] = 16'h0000;
	mel_filter_coefs[22][10] = 16'h0000;
	mel_filter_coefs[22][11] = 16'h0000;
	mel_filter_coefs[22][12] = 16'h0000;
	mel_filter_coefs[22][13] = 16'h0000;
	mel_filter_coefs[22][14] = 16'h0000;
	mel_filter_coefs[22][15] = 16'h0000;
	mel_filter_coefs[22][16] = 16'h0000;
	mel_filter_coefs[22][17] = 16'h0000;
	mel_filter_coefs[22][18] = 16'h0000;
	mel_filter_coefs[22][19] = 16'h0000;
	mel_filter_coefs[22][20] = 16'h0000;
	mel_filter_coefs[22][21] = 16'h0000;
	mel_filter_coefs[22][22] = 16'h0000;
	mel_filter_coefs[22][23] = 16'h0000;
	mel_filter_coefs[22][24] = 16'h0000;
	mel_filter_coefs[22][25] = 16'h0000;
	mel_filter_coefs[22][26] = 16'h0000;
	mel_filter_coefs[22][27] = 16'h0000;
	mel_filter_coefs[22][28] = 16'h0000;
	mel_filter_coefs[22][29] = 16'h0000;
	mel_filter_coefs[22][30] = 16'h0000;
	mel_filter_coefs[22][31] = 16'h0000;
	mel_filter_coefs[22][32] = 16'h0000;
	mel_filter_coefs[22][33] = 16'h0000;
	mel_filter_coefs[22][34] = 16'h0000;
	mel_filter_coefs[22][35] = 16'h0000;
	mel_filter_coefs[22][36] = 16'h0000;
	mel_filter_coefs[22][37] = 16'h0000;
	mel_filter_coefs[22][38] = 16'h0000;
	mel_filter_coefs[22][39] = 16'h0000;
	mel_filter_coefs[22][40] = 16'h0000;
	mel_filter_coefs[22][41] = 16'h0000;
	mel_filter_coefs[22][42] = 16'h0000;
	mel_filter_coefs[22][43] = 16'h0000;
	mel_filter_coefs[22][44] = 16'h0000;
	mel_filter_coefs[22][45] = 16'h0000;
	mel_filter_coefs[22][46] = 16'h0000;
	mel_filter_coefs[22][47] = 16'h0000;
	mel_filter_coefs[22][48] = 16'h0000;
	mel_filter_coefs[22][49] = 16'h0000;
	mel_filter_coefs[22][50] = 16'h0000;
	mel_filter_coefs[22][51] = 16'h0000;
	mel_filter_coefs[22][52] = 16'h0000;
	mel_filter_coefs[22][53] = 16'h0000;
	mel_filter_coefs[22][54] = 16'h0000;
	mel_filter_coefs[22][55] = 16'h0000;
	mel_filter_coefs[22][56] = 16'h0000;
	mel_filter_coefs[22][57] = 16'h0000;
	mel_filter_coefs[22][58] = 16'h0000;
	mel_filter_coefs[22][59] = 16'h0000;
	mel_filter_coefs[22][60] = 16'h0000;
	mel_filter_coefs[22][61] = 16'h0000;
	mel_filter_coefs[22][62] = 16'h0000;
	mel_filter_coefs[22][63] = 16'h0000;
	mel_filter_coefs[22][64] = 16'h0147;
	mel_filter_coefs[22][65] = 16'h18B0;
	mel_filter_coefs[22][66] = 16'h3019;
	mel_filter_coefs[22][67] = 16'h4781;
	mel_filter_coefs[22][68] = 16'h5EEA;
	mel_filter_coefs[22][69] = 16'h7653;
	mel_filter_coefs[22][70] = 16'h7316;
	mel_filter_coefs[22][71] = 16'h5D13;
	mel_filter_coefs[22][72] = 16'h470F;
	mel_filter_coefs[22][73] = 16'h310C;
	mel_filter_coefs[22][74] = 16'h1B08;
	mel_filter_coefs[22][75] = 16'h0505;
	mel_filter_coefs[22][76] = 16'h0000;
	mel_filter_coefs[22][77] = 16'h0000;
	mel_filter_coefs[22][78] = 16'h0000;
	mel_filter_coefs[22][79] = 16'h0000;
	mel_filter_coefs[22][80] = 16'h0000;
	mel_filter_coefs[22][81] = 16'h0000;
	mel_filter_coefs[22][82] = 16'h0000;
	mel_filter_coefs[22][83] = 16'h0000;
	mel_filter_coefs[22][84] = 16'h0000;
	mel_filter_coefs[22][85] = 16'h0000;
	mel_filter_coefs[22][86] = 16'h0000;
	mel_filter_coefs[22][87] = 16'h0000;
	mel_filter_coefs[22][88] = 16'h0000;
	mel_filter_coefs[22][89] = 16'h0000;
	mel_filter_coefs[22][90] = 16'h0000;
	mel_filter_coefs[22][91] = 16'h0000;
	mel_filter_coefs[22][92] = 16'h0000;
	mel_filter_coefs[22][93] = 16'h0000;
	mel_filter_coefs[22][94] = 16'h0000;
	mel_filter_coefs[22][95] = 16'h0000;
	mel_filter_coefs[22][96] = 16'h0000;
	mel_filter_coefs[22][97] = 16'h0000;
	mel_filter_coefs[22][98] = 16'h0000;
	mel_filter_coefs[22][99] = 16'h0000;
	mel_filter_coefs[22][100] = 16'h0000;
	mel_filter_coefs[22][101] = 16'h0000;
	mel_filter_coefs[22][102] = 16'h0000;
	mel_filter_coefs[22][103] = 16'h0000;
	mel_filter_coefs[22][104] = 16'h0000;
	mel_filter_coefs[22][105] = 16'h0000;
	mel_filter_coefs[22][106] = 16'h0000;
	mel_filter_coefs[22][107] = 16'h0000;
	mel_filter_coefs[22][108] = 16'h0000;
	mel_filter_coefs[22][109] = 16'h0000;
	mel_filter_coefs[22][110] = 16'h0000;
	mel_filter_coefs[22][111] = 16'h0000;
	mel_filter_coefs[22][112] = 16'h0000;
	mel_filter_coefs[22][113] = 16'h0000;
	mel_filter_coefs[22][114] = 16'h0000;
	mel_filter_coefs[22][115] = 16'h0000;
	mel_filter_coefs[22][116] = 16'h0000;
	mel_filter_coefs[22][117] = 16'h0000;
	mel_filter_coefs[22][118] = 16'h0000;
	mel_filter_coefs[22][119] = 16'h0000;
	mel_filter_coefs[22][120] = 16'h0000;
	mel_filter_coefs[22][121] = 16'h0000;
	mel_filter_coefs[22][122] = 16'h0000;
	mel_filter_coefs[22][123] = 16'h0000;
	mel_filter_coefs[22][124] = 16'h0000;
	mel_filter_coefs[22][125] = 16'h0000;
	mel_filter_coefs[22][126] = 16'h0000;
	mel_filter_coefs[22][127] = 16'h0000;
	mel_filter_coefs[22][128] = 16'h0000;
	mel_filter_coefs[22][129] = 16'h0000;
	mel_filter_coefs[22][130] = 16'h0000;
	mel_filter_coefs[22][131] = 16'h0000;
	mel_filter_coefs[22][132] = 16'h0000;
	mel_filter_coefs[22][133] = 16'h0000;
	mel_filter_coefs[22][134] = 16'h0000;
	mel_filter_coefs[22][135] = 16'h0000;
	mel_filter_coefs[22][136] = 16'h0000;
	mel_filter_coefs[22][137] = 16'h0000;
	mel_filter_coefs[22][138] = 16'h0000;
	mel_filter_coefs[22][139] = 16'h0000;
	mel_filter_coefs[22][140] = 16'h0000;
	mel_filter_coefs[22][141] = 16'h0000;
	mel_filter_coefs[22][142] = 16'h0000;
	mel_filter_coefs[22][143] = 16'h0000;
	mel_filter_coefs[22][144] = 16'h0000;
	mel_filter_coefs[22][145] = 16'h0000;
	mel_filter_coefs[22][146] = 16'h0000;
	mel_filter_coefs[22][147] = 16'h0000;
	mel_filter_coefs[22][148] = 16'h0000;
	mel_filter_coefs[22][149] = 16'h0000;
	mel_filter_coefs[22][150] = 16'h0000;
	mel_filter_coefs[22][151] = 16'h0000;
	mel_filter_coefs[22][152] = 16'h0000;
	mel_filter_coefs[22][153] = 16'h0000;
	mel_filter_coefs[22][154] = 16'h0000;
	mel_filter_coefs[22][155] = 16'h0000;
	mel_filter_coefs[22][156] = 16'h0000;
	mel_filter_coefs[22][157] = 16'h0000;
	mel_filter_coefs[22][158] = 16'h0000;
	mel_filter_coefs[22][159] = 16'h0000;
	mel_filter_coefs[22][160] = 16'h0000;
	mel_filter_coefs[22][161] = 16'h0000;
	mel_filter_coefs[22][162] = 16'h0000;
	mel_filter_coefs[22][163] = 16'h0000;
	mel_filter_coefs[22][164] = 16'h0000;
	mel_filter_coefs[22][165] = 16'h0000;
	mel_filter_coefs[22][166] = 16'h0000;
	mel_filter_coefs[22][167] = 16'h0000;
	mel_filter_coefs[22][168] = 16'h0000;
	mel_filter_coefs[22][169] = 16'h0000;
	mel_filter_coefs[22][170] = 16'h0000;
	mel_filter_coefs[22][171] = 16'h0000;
	mel_filter_coefs[22][172] = 16'h0000;
	mel_filter_coefs[22][173] = 16'h0000;
	mel_filter_coefs[22][174] = 16'h0000;
	mel_filter_coefs[22][175] = 16'h0000;
	mel_filter_coefs[22][176] = 16'h0000;
	mel_filter_coefs[22][177] = 16'h0000;
	mel_filter_coefs[22][178] = 16'h0000;
	mel_filter_coefs[22][179] = 16'h0000;
	mel_filter_coefs[22][180] = 16'h0000;
	mel_filter_coefs[22][181] = 16'h0000;
	mel_filter_coefs[22][182] = 16'h0000;
	mel_filter_coefs[22][183] = 16'h0000;
	mel_filter_coefs[22][184] = 16'h0000;
	mel_filter_coefs[22][185] = 16'h0000;
	mel_filter_coefs[22][186] = 16'h0000;
	mel_filter_coefs[22][187] = 16'h0000;
	mel_filter_coefs[22][188] = 16'h0000;
	mel_filter_coefs[22][189] = 16'h0000;
	mel_filter_coefs[22][190] = 16'h0000;
	mel_filter_coefs[22][191] = 16'h0000;
	mel_filter_coefs[22][192] = 16'h0000;
	mel_filter_coefs[22][193] = 16'h0000;
	mel_filter_coefs[22][194] = 16'h0000;
	mel_filter_coefs[22][195] = 16'h0000;
	mel_filter_coefs[22][196] = 16'h0000;
	mel_filter_coefs[22][197] = 16'h0000;
	mel_filter_coefs[22][198] = 16'h0000;
	mel_filter_coefs[22][199] = 16'h0000;
	mel_filter_coefs[22][200] = 16'h0000;
	mel_filter_coefs[22][201] = 16'h0000;
	mel_filter_coefs[22][202] = 16'h0000;
	mel_filter_coefs[22][203] = 16'h0000;
	mel_filter_coefs[22][204] = 16'h0000;
	mel_filter_coefs[22][205] = 16'h0000;
	mel_filter_coefs[22][206] = 16'h0000;
	mel_filter_coefs[22][207] = 16'h0000;
	mel_filter_coefs[22][208] = 16'h0000;
	mel_filter_coefs[22][209] = 16'h0000;
	mel_filter_coefs[22][210] = 16'h0000;
	mel_filter_coefs[22][211] = 16'h0000;
	mel_filter_coefs[22][212] = 16'h0000;
	mel_filter_coefs[22][213] = 16'h0000;
	mel_filter_coefs[22][214] = 16'h0000;
	mel_filter_coefs[22][215] = 16'h0000;
	mel_filter_coefs[22][216] = 16'h0000;
	mel_filter_coefs[22][217] = 16'h0000;
	mel_filter_coefs[22][218] = 16'h0000;
	mel_filter_coefs[22][219] = 16'h0000;
	mel_filter_coefs[22][220] = 16'h0000;
	mel_filter_coefs[22][221] = 16'h0000;
	mel_filter_coefs[22][222] = 16'h0000;
	mel_filter_coefs[22][223] = 16'h0000;
	mel_filter_coefs[22][224] = 16'h0000;
	mel_filter_coefs[22][225] = 16'h0000;
	mel_filter_coefs[22][226] = 16'h0000;
	mel_filter_coefs[22][227] = 16'h0000;
	mel_filter_coefs[22][228] = 16'h0000;
	mel_filter_coefs[22][229] = 16'h0000;
	mel_filter_coefs[22][230] = 16'h0000;
	mel_filter_coefs[22][231] = 16'h0000;
	mel_filter_coefs[22][232] = 16'h0000;
	mel_filter_coefs[22][233] = 16'h0000;
	mel_filter_coefs[22][234] = 16'h0000;
	mel_filter_coefs[22][235] = 16'h0000;
	mel_filter_coefs[22][236] = 16'h0000;
	mel_filter_coefs[22][237] = 16'h0000;
	mel_filter_coefs[22][238] = 16'h0000;
	mel_filter_coefs[22][239] = 16'h0000;
	mel_filter_coefs[22][240] = 16'h0000;
	mel_filter_coefs[22][241] = 16'h0000;
	mel_filter_coefs[22][242] = 16'h0000;
	mel_filter_coefs[22][243] = 16'h0000;
	mel_filter_coefs[22][244] = 16'h0000;
	mel_filter_coefs[22][245] = 16'h0000;
	mel_filter_coefs[22][246] = 16'h0000;
	mel_filter_coefs[22][247] = 16'h0000;
	mel_filter_coefs[22][248] = 16'h0000;
	mel_filter_coefs[22][249] = 16'h0000;
	mel_filter_coefs[22][250] = 16'h0000;
	mel_filter_coefs[22][251] = 16'h0000;
	mel_filter_coefs[22][252] = 16'h0000;
	mel_filter_coefs[22][253] = 16'h0000;
	mel_filter_coefs[22][254] = 16'h0000;
	mel_filter_coefs[22][255] = 16'h0000;
	mel_filter_coefs[23][0] = 16'h0000;
	mel_filter_coefs[23][1] = 16'h0000;
	mel_filter_coefs[23][2] = 16'h0000;
	mel_filter_coefs[23][3] = 16'h0000;
	mel_filter_coefs[23][4] = 16'h0000;
	mel_filter_coefs[23][5] = 16'h0000;
	mel_filter_coefs[23][6] = 16'h0000;
	mel_filter_coefs[23][7] = 16'h0000;
	mel_filter_coefs[23][8] = 16'h0000;
	mel_filter_coefs[23][9] = 16'h0000;
	mel_filter_coefs[23][10] = 16'h0000;
	mel_filter_coefs[23][11] = 16'h0000;
	mel_filter_coefs[23][12] = 16'h0000;
	mel_filter_coefs[23][13] = 16'h0000;
	mel_filter_coefs[23][14] = 16'h0000;
	mel_filter_coefs[23][15] = 16'h0000;
	mel_filter_coefs[23][16] = 16'h0000;
	mel_filter_coefs[23][17] = 16'h0000;
	mel_filter_coefs[23][18] = 16'h0000;
	mel_filter_coefs[23][19] = 16'h0000;
	mel_filter_coefs[23][20] = 16'h0000;
	mel_filter_coefs[23][21] = 16'h0000;
	mel_filter_coefs[23][22] = 16'h0000;
	mel_filter_coefs[23][23] = 16'h0000;
	mel_filter_coefs[23][24] = 16'h0000;
	mel_filter_coefs[23][25] = 16'h0000;
	mel_filter_coefs[23][26] = 16'h0000;
	mel_filter_coefs[23][27] = 16'h0000;
	mel_filter_coefs[23][28] = 16'h0000;
	mel_filter_coefs[23][29] = 16'h0000;
	mel_filter_coefs[23][30] = 16'h0000;
	mel_filter_coefs[23][31] = 16'h0000;
	mel_filter_coefs[23][32] = 16'h0000;
	mel_filter_coefs[23][33] = 16'h0000;
	mel_filter_coefs[23][34] = 16'h0000;
	mel_filter_coefs[23][35] = 16'h0000;
	mel_filter_coefs[23][36] = 16'h0000;
	mel_filter_coefs[23][37] = 16'h0000;
	mel_filter_coefs[23][38] = 16'h0000;
	mel_filter_coefs[23][39] = 16'h0000;
	mel_filter_coefs[23][40] = 16'h0000;
	mel_filter_coefs[23][41] = 16'h0000;
	mel_filter_coefs[23][42] = 16'h0000;
	mel_filter_coefs[23][43] = 16'h0000;
	mel_filter_coefs[23][44] = 16'h0000;
	mel_filter_coefs[23][45] = 16'h0000;
	mel_filter_coefs[23][46] = 16'h0000;
	mel_filter_coefs[23][47] = 16'h0000;
	mel_filter_coefs[23][48] = 16'h0000;
	mel_filter_coefs[23][49] = 16'h0000;
	mel_filter_coefs[23][50] = 16'h0000;
	mel_filter_coefs[23][51] = 16'h0000;
	mel_filter_coefs[23][52] = 16'h0000;
	mel_filter_coefs[23][53] = 16'h0000;
	mel_filter_coefs[23][54] = 16'h0000;
	mel_filter_coefs[23][55] = 16'h0000;
	mel_filter_coefs[23][56] = 16'h0000;
	mel_filter_coefs[23][57] = 16'h0000;
	mel_filter_coefs[23][58] = 16'h0000;
	mel_filter_coefs[23][59] = 16'h0000;
	mel_filter_coefs[23][60] = 16'h0000;
	mel_filter_coefs[23][61] = 16'h0000;
	mel_filter_coefs[23][62] = 16'h0000;
	mel_filter_coefs[23][63] = 16'h0000;
	mel_filter_coefs[23][64] = 16'h0000;
	mel_filter_coefs[23][65] = 16'h0000;
	mel_filter_coefs[23][66] = 16'h0000;
	mel_filter_coefs[23][67] = 16'h0000;
	mel_filter_coefs[23][68] = 16'h0000;
	mel_filter_coefs[23][69] = 16'h0000;
	mel_filter_coefs[23][70] = 16'h0CEA;
	mel_filter_coefs[23][71] = 16'h22ED;
	mel_filter_coefs[23][72] = 16'h38F1;
	mel_filter_coefs[23][73] = 16'h4EF4;
	mel_filter_coefs[23][74] = 16'h64F8;
	mel_filter_coefs[23][75] = 16'h7AFB;
	mel_filter_coefs[23][76] = 16'h7005;
	mel_filter_coefs[23][77] = 16'h5B51;
	mel_filter_coefs[23][78] = 16'h469E;
	mel_filter_coefs[23][79] = 16'h31EA;
	mel_filter_coefs[23][80] = 16'h1D37;
	mel_filter_coefs[23][81] = 16'h0883;
	mel_filter_coefs[23][82] = 16'h0000;
	mel_filter_coefs[23][83] = 16'h0000;
	mel_filter_coefs[23][84] = 16'h0000;
	mel_filter_coefs[23][85] = 16'h0000;
	mel_filter_coefs[23][86] = 16'h0000;
	mel_filter_coefs[23][87] = 16'h0000;
	mel_filter_coefs[23][88] = 16'h0000;
	mel_filter_coefs[23][89] = 16'h0000;
	mel_filter_coefs[23][90] = 16'h0000;
	mel_filter_coefs[23][91] = 16'h0000;
	mel_filter_coefs[23][92] = 16'h0000;
	mel_filter_coefs[23][93] = 16'h0000;
	mel_filter_coefs[23][94] = 16'h0000;
	mel_filter_coefs[23][95] = 16'h0000;
	mel_filter_coefs[23][96] = 16'h0000;
	mel_filter_coefs[23][97] = 16'h0000;
	mel_filter_coefs[23][98] = 16'h0000;
	mel_filter_coefs[23][99] = 16'h0000;
	mel_filter_coefs[23][100] = 16'h0000;
	mel_filter_coefs[23][101] = 16'h0000;
	mel_filter_coefs[23][102] = 16'h0000;
	mel_filter_coefs[23][103] = 16'h0000;
	mel_filter_coefs[23][104] = 16'h0000;
	mel_filter_coefs[23][105] = 16'h0000;
	mel_filter_coefs[23][106] = 16'h0000;
	mel_filter_coefs[23][107] = 16'h0000;
	mel_filter_coefs[23][108] = 16'h0000;
	mel_filter_coefs[23][109] = 16'h0000;
	mel_filter_coefs[23][110] = 16'h0000;
	mel_filter_coefs[23][111] = 16'h0000;
	mel_filter_coefs[23][112] = 16'h0000;
	mel_filter_coefs[23][113] = 16'h0000;
	mel_filter_coefs[23][114] = 16'h0000;
	mel_filter_coefs[23][115] = 16'h0000;
	mel_filter_coefs[23][116] = 16'h0000;
	mel_filter_coefs[23][117] = 16'h0000;
	mel_filter_coefs[23][118] = 16'h0000;
	mel_filter_coefs[23][119] = 16'h0000;
	mel_filter_coefs[23][120] = 16'h0000;
	mel_filter_coefs[23][121] = 16'h0000;
	mel_filter_coefs[23][122] = 16'h0000;
	mel_filter_coefs[23][123] = 16'h0000;
	mel_filter_coefs[23][124] = 16'h0000;
	mel_filter_coefs[23][125] = 16'h0000;
	mel_filter_coefs[23][126] = 16'h0000;
	mel_filter_coefs[23][127] = 16'h0000;
	mel_filter_coefs[23][128] = 16'h0000;
	mel_filter_coefs[23][129] = 16'h0000;
	mel_filter_coefs[23][130] = 16'h0000;
	mel_filter_coefs[23][131] = 16'h0000;
	mel_filter_coefs[23][132] = 16'h0000;
	mel_filter_coefs[23][133] = 16'h0000;
	mel_filter_coefs[23][134] = 16'h0000;
	mel_filter_coefs[23][135] = 16'h0000;
	mel_filter_coefs[23][136] = 16'h0000;
	mel_filter_coefs[23][137] = 16'h0000;
	mel_filter_coefs[23][138] = 16'h0000;
	mel_filter_coefs[23][139] = 16'h0000;
	mel_filter_coefs[23][140] = 16'h0000;
	mel_filter_coefs[23][141] = 16'h0000;
	mel_filter_coefs[23][142] = 16'h0000;
	mel_filter_coefs[23][143] = 16'h0000;
	mel_filter_coefs[23][144] = 16'h0000;
	mel_filter_coefs[23][145] = 16'h0000;
	mel_filter_coefs[23][146] = 16'h0000;
	mel_filter_coefs[23][147] = 16'h0000;
	mel_filter_coefs[23][148] = 16'h0000;
	mel_filter_coefs[23][149] = 16'h0000;
	mel_filter_coefs[23][150] = 16'h0000;
	mel_filter_coefs[23][151] = 16'h0000;
	mel_filter_coefs[23][152] = 16'h0000;
	mel_filter_coefs[23][153] = 16'h0000;
	mel_filter_coefs[23][154] = 16'h0000;
	mel_filter_coefs[23][155] = 16'h0000;
	mel_filter_coefs[23][156] = 16'h0000;
	mel_filter_coefs[23][157] = 16'h0000;
	mel_filter_coefs[23][158] = 16'h0000;
	mel_filter_coefs[23][159] = 16'h0000;
	mel_filter_coefs[23][160] = 16'h0000;
	mel_filter_coefs[23][161] = 16'h0000;
	mel_filter_coefs[23][162] = 16'h0000;
	mel_filter_coefs[23][163] = 16'h0000;
	mel_filter_coefs[23][164] = 16'h0000;
	mel_filter_coefs[23][165] = 16'h0000;
	mel_filter_coefs[23][166] = 16'h0000;
	mel_filter_coefs[23][167] = 16'h0000;
	mel_filter_coefs[23][168] = 16'h0000;
	mel_filter_coefs[23][169] = 16'h0000;
	mel_filter_coefs[23][170] = 16'h0000;
	mel_filter_coefs[23][171] = 16'h0000;
	mel_filter_coefs[23][172] = 16'h0000;
	mel_filter_coefs[23][173] = 16'h0000;
	mel_filter_coefs[23][174] = 16'h0000;
	mel_filter_coefs[23][175] = 16'h0000;
	mel_filter_coefs[23][176] = 16'h0000;
	mel_filter_coefs[23][177] = 16'h0000;
	mel_filter_coefs[23][178] = 16'h0000;
	mel_filter_coefs[23][179] = 16'h0000;
	mel_filter_coefs[23][180] = 16'h0000;
	mel_filter_coefs[23][181] = 16'h0000;
	mel_filter_coefs[23][182] = 16'h0000;
	mel_filter_coefs[23][183] = 16'h0000;
	mel_filter_coefs[23][184] = 16'h0000;
	mel_filter_coefs[23][185] = 16'h0000;
	mel_filter_coefs[23][186] = 16'h0000;
	mel_filter_coefs[23][187] = 16'h0000;
	mel_filter_coefs[23][188] = 16'h0000;
	mel_filter_coefs[23][189] = 16'h0000;
	mel_filter_coefs[23][190] = 16'h0000;
	mel_filter_coefs[23][191] = 16'h0000;
	mel_filter_coefs[23][192] = 16'h0000;
	mel_filter_coefs[23][193] = 16'h0000;
	mel_filter_coefs[23][194] = 16'h0000;
	mel_filter_coefs[23][195] = 16'h0000;
	mel_filter_coefs[23][196] = 16'h0000;
	mel_filter_coefs[23][197] = 16'h0000;
	mel_filter_coefs[23][198] = 16'h0000;
	mel_filter_coefs[23][199] = 16'h0000;
	mel_filter_coefs[23][200] = 16'h0000;
	mel_filter_coefs[23][201] = 16'h0000;
	mel_filter_coefs[23][202] = 16'h0000;
	mel_filter_coefs[23][203] = 16'h0000;
	mel_filter_coefs[23][204] = 16'h0000;
	mel_filter_coefs[23][205] = 16'h0000;
	mel_filter_coefs[23][206] = 16'h0000;
	mel_filter_coefs[23][207] = 16'h0000;
	mel_filter_coefs[23][208] = 16'h0000;
	mel_filter_coefs[23][209] = 16'h0000;
	mel_filter_coefs[23][210] = 16'h0000;
	mel_filter_coefs[23][211] = 16'h0000;
	mel_filter_coefs[23][212] = 16'h0000;
	mel_filter_coefs[23][213] = 16'h0000;
	mel_filter_coefs[23][214] = 16'h0000;
	mel_filter_coefs[23][215] = 16'h0000;
	mel_filter_coefs[23][216] = 16'h0000;
	mel_filter_coefs[23][217] = 16'h0000;
	mel_filter_coefs[23][218] = 16'h0000;
	mel_filter_coefs[23][219] = 16'h0000;
	mel_filter_coefs[23][220] = 16'h0000;
	mel_filter_coefs[23][221] = 16'h0000;
	mel_filter_coefs[23][222] = 16'h0000;
	mel_filter_coefs[23][223] = 16'h0000;
	mel_filter_coefs[23][224] = 16'h0000;
	mel_filter_coefs[23][225] = 16'h0000;
	mel_filter_coefs[23][226] = 16'h0000;
	mel_filter_coefs[23][227] = 16'h0000;
	mel_filter_coefs[23][228] = 16'h0000;
	mel_filter_coefs[23][229] = 16'h0000;
	mel_filter_coefs[23][230] = 16'h0000;
	mel_filter_coefs[23][231] = 16'h0000;
	mel_filter_coefs[23][232] = 16'h0000;
	mel_filter_coefs[23][233] = 16'h0000;
	mel_filter_coefs[23][234] = 16'h0000;
	mel_filter_coefs[23][235] = 16'h0000;
	mel_filter_coefs[23][236] = 16'h0000;
	mel_filter_coefs[23][237] = 16'h0000;
	mel_filter_coefs[23][238] = 16'h0000;
	mel_filter_coefs[23][239] = 16'h0000;
	mel_filter_coefs[23][240] = 16'h0000;
	mel_filter_coefs[23][241] = 16'h0000;
	mel_filter_coefs[23][242] = 16'h0000;
	mel_filter_coefs[23][243] = 16'h0000;
	mel_filter_coefs[23][244] = 16'h0000;
	mel_filter_coefs[23][245] = 16'h0000;
	mel_filter_coefs[23][246] = 16'h0000;
	mel_filter_coefs[23][247] = 16'h0000;
	mel_filter_coefs[23][248] = 16'h0000;
	mel_filter_coefs[23][249] = 16'h0000;
	mel_filter_coefs[23][250] = 16'h0000;
	mel_filter_coefs[23][251] = 16'h0000;
	mel_filter_coefs[23][252] = 16'h0000;
	mel_filter_coefs[23][253] = 16'h0000;
	mel_filter_coefs[23][254] = 16'h0000;
	mel_filter_coefs[23][255] = 16'h0000;
	mel_filter_coefs[24][0] = 16'h0000;
	mel_filter_coefs[24][1] = 16'h0000;
	mel_filter_coefs[24][2] = 16'h0000;
	mel_filter_coefs[24][3] = 16'h0000;
	mel_filter_coefs[24][4] = 16'h0000;
	mel_filter_coefs[24][5] = 16'h0000;
	mel_filter_coefs[24][6] = 16'h0000;
	mel_filter_coefs[24][7] = 16'h0000;
	mel_filter_coefs[24][8] = 16'h0000;
	mel_filter_coefs[24][9] = 16'h0000;
	mel_filter_coefs[24][10] = 16'h0000;
	mel_filter_coefs[24][11] = 16'h0000;
	mel_filter_coefs[24][12] = 16'h0000;
	mel_filter_coefs[24][13] = 16'h0000;
	mel_filter_coefs[24][14] = 16'h0000;
	mel_filter_coefs[24][15] = 16'h0000;
	mel_filter_coefs[24][16] = 16'h0000;
	mel_filter_coefs[24][17] = 16'h0000;
	mel_filter_coefs[24][18] = 16'h0000;
	mel_filter_coefs[24][19] = 16'h0000;
	mel_filter_coefs[24][20] = 16'h0000;
	mel_filter_coefs[24][21] = 16'h0000;
	mel_filter_coefs[24][22] = 16'h0000;
	mel_filter_coefs[24][23] = 16'h0000;
	mel_filter_coefs[24][24] = 16'h0000;
	mel_filter_coefs[24][25] = 16'h0000;
	mel_filter_coefs[24][26] = 16'h0000;
	mel_filter_coefs[24][27] = 16'h0000;
	mel_filter_coefs[24][28] = 16'h0000;
	mel_filter_coefs[24][29] = 16'h0000;
	mel_filter_coefs[24][30] = 16'h0000;
	mel_filter_coefs[24][31] = 16'h0000;
	mel_filter_coefs[24][32] = 16'h0000;
	mel_filter_coefs[24][33] = 16'h0000;
	mel_filter_coefs[24][34] = 16'h0000;
	mel_filter_coefs[24][35] = 16'h0000;
	mel_filter_coefs[24][36] = 16'h0000;
	mel_filter_coefs[24][37] = 16'h0000;
	mel_filter_coefs[24][38] = 16'h0000;
	mel_filter_coefs[24][39] = 16'h0000;
	mel_filter_coefs[24][40] = 16'h0000;
	mel_filter_coefs[24][41] = 16'h0000;
	mel_filter_coefs[24][42] = 16'h0000;
	mel_filter_coefs[24][43] = 16'h0000;
	mel_filter_coefs[24][44] = 16'h0000;
	mel_filter_coefs[24][45] = 16'h0000;
	mel_filter_coefs[24][46] = 16'h0000;
	mel_filter_coefs[24][47] = 16'h0000;
	mel_filter_coefs[24][48] = 16'h0000;
	mel_filter_coefs[24][49] = 16'h0000;
	mel_filter_coefs[24][50] = 16'h0000;
	mel_filter_coefs[24][51] = 16'h0000;
	mel_filter_coefs[24][52] = 16'h0000;
	mel_filter_coefs[24][53] = 16'h0000;
	mel_filter_coefs[24][54] = 16'h0000;
	mel_filter_coefs[24][55] = 16'h0000;
	mel_filter_coefs[24][56] = 16'h0000;
	mel_filter_coefs[24][57] = 16'h0000;
	mel_filter_coefs[24][58] = 16'h0000;
	mel_filter_coefs[24][59] = 16'h0000;
	mel_filter_coefs[24][60] = 16'h0000;
	mel_filter_coefs[24][61] = 16'h0000;
	mel_filter_coefs[24][62] = 16'h0000;
	mel_filter_coefs[24][63] = 16'h0000;
	mel_filter_coefs[24][64] = 16'h0000;
	mel_filter_coefs[24][65] = 16'h0000;
	mel_filter_coefs[24][66] = 16'h0000;
	mel_filter_coefs[24][67] = 16'h0000;
	mel_filter_coefs[24][68] = 16'h0000;
	mel_filter_coefs[24][69] = 16'h0000;
	mel_filter_coefs[24][70] = 16'h0000;
	mel_filter_coefs[24][71] = 16'h0000;
	mel_filter_coefs[24][72] = 16'h0000;
	mel_filter_coefs[24][73] = 16'h0000;
	mel_filter_coefs[24][74] = 16'h0000;
	mel_filter_coefs[24][75] = 16'h0000;
	mel_filter_coefs[24][76] = 16'h0FFB;
	mel_filter_coefs[24][77] = 16'h24AF;
	mel_filter_coefs[24][78] = 16'h3962;
	mel_filter_coefs[24][79] = 16'h4E16;
	mel_filter_coefs[24][80] = 16'h62C9;
	mel_filter_coefs[24][81] = 16'h777D;
	mel_filter_coefs[24][82] = 16'h748A;
	mel_filter_coefs[24][83] = 16'h6112;
	mel_filter_coefs[24][84] = 16'h4D9B;
	mel_filter_coefs[24][85] = 16'h3A23;
	mel_filter_coefs[24][86] = 16'h26AC;
	mel_filter_coefs[24][87] = 16'h1334;
	mel_filter_coefs[24][88] = 16'h0000;
	mel_filter_coefs[24][89] = 16'h0000;
	mel_filter_coefs[24][90] = 16'h0000;
	mel_filter_coefs[24][91] = 16'h0000;
	mel_filter_coefs[24][92] = 16'h0000;
	mel_filter_coefs[24][93] = 16'h0000;
	mel_filter_coefs[24][94] = 16'h0000;
	mel_filter_coefs[24][95] = 16'h0000;
	mel_filter_coefs[24][96] = 16'h0000;
	mel_filter_coefs[24][97] = 16'h0000;
	mel_filter_coefs[24][98] = 16'h0000;
	mel_filter_coefs[24][99] = 16'h0000;
	mel_filter_coefs[24][100] = 16'h0000;
	mel_filter_coefs[24][101] = 16'h0000;
	mel_filter_coefs[24][102] = 16'h0000;
	mel_filter_coefs[24][103] = 16'h0000;
	mel_filter_coefs[24][104] = 16'h0000;
	mel_filter_coefs[24][105] = 16'h0000;
	mel_filter_coefs[24][106] = 16'h0000;
	mel_filter_coefs[24][107] = 16'h0000;
	mel_filter_coefs[24][108] = 16'h0000;
	mel_filter_coefs[24][109] = 16'h0000;
	mel_filter_coefs[24][110] = 16'h0000;
	mel_filter_coefs[24][111] = 16'h0000;
	mel_filter_coefs[24][112] = 16'h0000;
	mel_filter_coefs[24][113] = 16'h0000;
	mel_filter_coefs[24][114] = 16'h0000;
	mel_filter_coefs[24][115] = 16'h0000;
	mel_filter_coefs[24][116] = 16'h0000;
	mel_filter_coefs[24][117] = 16'h0000;
	mel_filter_coefs[24][118] = 16'h0000;
	mel_filter_coefs[24][119] = 16'h0000;
	mel_filter_coefs[24][120] = 16'h0000;
	mel_filter_coefs[24][121] = 16'h0000;
	mel_filter_coefs[24][122] = 16'h0000;
	mel_filter_coefs[24][123] = 16'h0000;
	mel_filter_coefs[24][124] = 16'h0000;
	mel_filter_coefs[24][125] = 16'h0000;
	mel_filter_coefs[24][126] = 16'h0000;
	mel_filter_coefs[24][127] = 16'h0000;
	mel_filter_coefs[24][128] = 16'h0000;
	mel_filter_coefs[24][129] = 16'h0000;
	mel_filter_coefs[24][130] = 16'h0000;
	mel_filter_coefs[24][131] = 16'h0000;
	mel_filter_coefs[24][132] = 16'h0000;
	mel_filter_coefs[24][133] = 16'h0000;
	mel_filter_coefs[24][134] = 16'h0000;
	mel_filter_coefs[24][135] = 16'h0000;
	mel_filter_coefs[24][136] = 16'h0000;
	mel_filter_coefs[24][137] = 16'h0000;
	mel_filter_coefs[24][138] = 16'h0000;
	mel_filter_coefs[24][139] = 16'h0000;
	mel_filter_coefs[24][140] = 16'h0000;
	mel_filter_coefs[24][141] = 16'h0000;
	mel_filter_coefs[24][142] = 16'h0000;
	mel_filter_coefs[24][143] = 16'h0000;
	mel_filter_coefs[24][144] = 16'h0000;
	mel_filter_coefs[24][145] = 16'h0000;
	mel_filter_coefs[24][146] = 16'h0000;
	mel_filter_coefs[24][147] = 16'h0000;
	mel_filter_coefs[24][148] = 16'h0000;
	mel_filter_coefs[24][149] = 16'h0000;
	mel_filter_coefs[24][150] = 16'h0000;
	mel_filter_coefs[24][151] = 16'h0000;
	mel_filter_coefs[24][152] = 16'h0000;
	mel_filter_coefs[24][153] = 16'h0000;
	mel_filter_coefs[24][154] = 16'h0000;
	mel_filter_coefs[24][155] = 16'h0000;
	mel_filter_coefs[24][156] = 16'h0000;
	mel_filter_coefs[24][157] = 16'h0000;
	mel_filter_coefs[24][158] = 16'h0000;
	mel_filter_coefs[24][159] = 16'h0000;
	mel_filter_coefs[24][160] = 16'h0000;
	mel_filter_coefs[24][161] = 16'h0000;
	mel_filter_coefs[24][162] = 16'h0000;
	mel_filter_coefs[24][163] = 16'h0000;
	mel_filter_coefs[24][164] = 16'h0000;
	mel_filter_coefs[24][165] = 16'h0000;
	mel_filter_coefs[24][166] = 16'h0000;
	mel_filter_coefs[24][167] = 16'h0000;
	mel_filter_coefs[24][168] = 16'h0000;
	mel_filter_coefs[24][169] = 16'h0000;
	mel_filter_coefs[24][170] = 16'h0000;
	mel_filter_coefs[24][171] = 16'h0000;
	mel_filter_coefs[24][172] = 16'h0000;
	mel_filter_coefs[24][173] = 16'h0000;
	mel_filter_coefs[24][174] = 16'h0000;
	mel_filter_coefs[24][175] = 16'h0000;
	mel_filter_coefs[24][176] = 16'h0000;
	mel_filter_coefs[24][177] = 16'h0000;
	mel_filter_coefs[24][178] = 16'h0000;
	mel_filter_coefs[24][179] = 16'h0000;
	mel_filter_coefs[24][180] = 16'h0000;
	mel_filter_coefs[24][181] = 16'h0000;
	mel_filter_coefs[24][182] = 16'h0000;
	mel_filter_coefs[24][183] = 16'h0000;
	mel_filter_coefs[24][184] = 16'h0000;
	mel_filter_coefs[24][185] = 16'h0000;
	mel_filter_coefs[24][186] = 16'h0000;
	mel_filter_coefs[24][187] = 16'h0000;
	mel_filter_coefs[24][188] = 16'h0000;
	mel_filter_coefs[24][189] = 16'h0000;
	mel_filter_coefs[24][190] = 16'h0000;
	mel_filter_coefs[24][191] = 16'h0000;
	mel_filter_coefs[24][192] = 16'h0000;
	mel_filter_coefs[24][193] = 16'h0000;
	mel_filter_coefs[24][194] = 16'h0000;
	mel_filter_coefs[24][195] = 16'h0000;
	mel_filter_coefs[24][196] = 16'h0000;
	mel_filter_coefs[24][197] = 16'h0000;
	mel_filter_coefs[24][198] = 16'h0000;
	mel_filter_coefs[24][199] = 16'h0000;
	mel_filter_coefs[24][200] = 16'h0000;
	mel_filter_coefs[24][201] = 16'h0000;
	mel_filter_coefs[24][202] = 16'h0000;
	mel_filter_coefs[24][203] = 16'h0000;
	mel_filter_coefs[24][204] = 16'h0000;
	mel_filter_coefs[24][205] = 16'h0000;
	mel_filter_coefs[24][206] = 16'h0000;
	mel_filter_coefs[24][207] = 16'h0000;
	mel_filter_coefs[24][208] = 16'h0000;
	mel_filter_coefs[24][209] = 16'h0000;
	mel_filter_coefs[24][210] = 16'h0000;
	mel_filter_coefs[24][211] = 16'h0000;
	mel_filter_coefs[24][212] = 16'h0000;
	mel_filter_coefs[24][213] = 16'h0000;
	mel_filter_coefs[24][214] = 16'h0000;
	mel_filter_coefs[24][215] = 16'h0000;
	mel_filter_coefs[24][216] = 16'h0000;
	mel_filter_coefs[24][217] = 16'h0000;
	mel_filter_coefs[24][218] = 16'h0000;
	mel_filter_coefs[24][219] = 16'h0000;
	mel_filter_coefs[24][220] = 16'h0000;
	mel_filter_coefs[24][221] = 16'h0000;
	mel_filter_coefs[24][222] = 16'h0000;
	mel_filter_coefs[24][223] = 16'h0000;
	mel_filter_coefs[24][224] = 16'h0000;
	mel_filter_coefs[24][225] = 16'h0000;
	mel_filter_coefs[24][226] = 16'h0000;
	mel_filter_coefs[24][227] = 16'h0000;
	mel_filter_coefs[24][228] = 16'h0000;
	mel_filter_coefs[24][229] = 16'h0000;
	mel_filter_coefs[24][230] = 16'h0000;
	mel_filter_coefs[24][231] = 16'h0000;
	mel_filter_coefs[24][232] = 16'h0000;
	mel_filter_coefs[24][233] = 16'h0000;
	mel_filter_coefs[24][234] = 16'h0000;
	mel_filter_coefs[24][235] = 16'h0000;
	mel_filter_coefs[24][236] = 16'h0000;
	mel_filter_coefs[24][237] = 16'h0000;
	mel_filter_coefs[24][238] = 16'h0000;
	mel_filter_coefs[24][239] = 16'h0000;
	mel_filter_coefs[24][240] = 16'h0000;
	mel_filter_coefs[24][241] = 16'h0000;
	mel_filter_coefs[24][242] = 16'h0000;
	mel_filter_coefs[24][243] = 16'h0000;
	mel_filter_coefs[24][244] = 16'h0000;
	mel_filter_coefs[24][245] = 16'h0000;
	mel_filter_coefs[24][246] = 16'h0000;
	mel_filter_coefs[24][247] = 16'h0000;
	mel_filter_coefs[24][248] = 16'h0000;
	mel_filter_coefs[24][249] = 16'h0000;
	mel_filter_coefs[24][250] = 16'h0000;
	mel_filter_coefs[24][251] = 16'h0000;
	mel_filter_coefs[24][252] = 16'h0000;
	mel_filter_coefs[24][253] = 16'h0000;
	mel_filter_coefs[24][254] = 16'h0000;
	mel_filter_coefs[24][255] = 16'h0000;
	mel_filter_coefs[25][0] = 16'h0000;
	mel_filter_coefs[25][1] = 16'h0000;
	mel_filter_coefs[25][2] = 16'h0000;
	mel_filter_coefs[25][3] = 16'h0000;
	mel_filter_coefs[25][4] = 16'h0000;
	mel_filter_coefs[25][5] = 16'h0000;
	mel_filter_coefs[25][6] = 16'h0000;
	mel_filter_coefs[25][7] = 16'h0000;
	mel_filter_coefs[25][8] = 16'h0000;
	mel_filter_coefs[25][9] = 16'h0000;
	mel_filter_coefs[25][10] = 16'h0000;
	mel_filter_coefs[25][11] = 16'h0000;
	mel_filter_coefs[25][12] = 16'h0000;
	mel_filter_coefs[25][13] = 16'h0000;
	mel_filter_coefs[25][14] = 16'h0000;
	mel_filter_coefs[25][15] = 16'h0000;
	mel_filter_coefs[25][16] = 16'h0000;
	mel_filter_coefs[25][17] = 16'h0000;
	mel_filter_coefs[25][18] = 16'h0000;
	mel_filter_coefs[25][19] = 16'h0000;
	mel_filter_coefs[25][20] = 16'h0000;
	mel_filter_coefs[25][21] = 16'h0000;
	mel_filter_coefs[25][22] = 16'h0000;
	mel_filter_coefs[25][23] = 16'h0000;
	mel_filter_coefs[25][24] = 16'h0000;
	mel_filter_coefs[25][25] = 16'h0000;
	mel_filter_coefs[25][26] = 16'h0000;
	mel_filter_coefs[25][27] = 16'h0000;
	mel_filter_coefs[25][28] = 16'h0000;
	mel_filter_coefs[25][29] = 16'h0000;
	mel_filter_coefs[25][30] = 16'h0000;
	mel_filter_coefs[25][31] = 16'h0000;
	mel_filter_coefs[25][32] = 16'h0000;
	mel_filter_coefs[25][33] = 16'h0000;
	mel_filter_coefs[25][34] = 16'h0000;
	mel_filter_coefs[25][35] = 16'h0000;
	mel_filter_coefs[25][36] = 16'h0000;
	mel_filter_coefs[25][37] = 16'h0000;
	mel_filter_coefs[25][38] = 16'h0000;
	mel_filter_coefs[25][39] = 16'h0000;
	mel_filter_coefs[25][40] = 16'h0000;
	mel_filter_coefs[25][41] = 16'h0000;
	mel_filter_coefs[25][42] = 16'h0000;
	mel_filter_coefs[25][43] = 16'h0000;
	mel_filter_coefs[25][44] = 16'h0000;
	mel_filter_coefs[25][45] = 16'h0000;
	mel_filter_coefs[25][46] = 16'h0000;
	mel_filter_coefs[25][47] = 16'h0000;
	mel_filter_coefs[25][48] = 16'h0000;
	mel_filter_coefs[25][49] = 16'h0000;
	mel_filter_coefs[25][50] = 16'h0000;
	mel_filter_coefs[25][51] = 16'h0000;
	mel_filter_coefs[25][52] = 16'h0000;
	mel_filter_coefs[25][53] = 16'h0000;
	mel_filter_coefs[25][54] = 16'h0000;
	mel_filter_coefs[25][55] = 16'h0000;
	mel_filter_coefs[25][56] = 16'h0000;
	mel_filter_coefs[25][57] = 16'h0000;
	mel_filter_coefs[25][58] = 16'h0000;
	mel_filter_coefs[25][59] = 16'h0000;
	mel_filter_coefs[25][60] = 16'h0000;
	mel_filter_coefs[25][61] = 16'h0000;
	mel_filter_coefs[25][62] = 16'h0000;
	mel_filter_coefs[25][63] = 16'h0000;
	mel_filter_coefs[25][64] = 16'h0000;
	mel_filter_coefs[25][65] = 16'h0000;
	mel_filter_coefs[25][66] = 16'h0000;
	mel_filter_coefs[25][67] = 16'h0000;
	mel_filter_coefs[25][68] = 16'h0000;
	mel_filter_coefs[25][69] = 16'h0000;
	mel_filter_coefs[25][70] = 16'h0000;
	mel_filter_coefs[25][71] = 16'h0000;
	mel_filter_coefs[25][72] = 16'h0000;
	mel_filter_coefs[25][73] = 16'h0000;
	mel_filter_coefs[25][74] = 16'h0000;
	mel_filter_coefs[25][75] = 16'h0000;
	mel_filter_coefs[25][76] = 16'h0000;
	mel_filter_coefs[25][77] = 16'h0000;
	mel_filter_coefs[25][78] = 16'h0000;
	mel_filter_coefs[25][79] = 16'h0000;
	mel_filter_coefs[25][80] = 16'h0000;
	mel_filter_coefs[25][81] = 16'h0000;
	mel_filter_coefs[25][82] = 16'h0B76;
	mel_filter_coefs[25][83] = 16'h1EEE;
	mel_filter_coefs[25][84] = 16'h3265;
	mel_filter_coefs[25][85] = 16'h45DD;
	mel_filter_coefs[25][86] = 16'h5954;
	mel_filter_coefs[25][87] = 16'h6CCC;
	mel_filter_coefs[25][88] = 16'h7FC1;
	mel_filter_coefs[25][89] = 16'h6D72;
	mel_filter_coefs[25][90] = 16'h5B24;
	mel_filter_coefs[25][91] = 16'h48D5;
	mel_filter_coefs[25][92] = 16'h3687;
	mel_filter_coefs[25][93] = 16'h2438;
	mel_filter_coefs[25][94] = 16'h11EA;
	mel_filter_coefs[25][95] = 16'h0000;
	mel_filter_coefs[25][96] = 16'h0000;
	mel_filter_coefs[25][97] = 16'h0000;
	mel_filter_coefs[25][98] = 16'h0000;
	mel_filter_coefs[25][99] = 16'h0000;
	mel_filter_coefs[25][100] = 16'h0000;
	mel_filter_coefs[25][101] = 16'h0000;
	mel_filter_coefs[25][102] = 16'h0000;
	mel_filter_coefs[25][103] = 16'h0000;
	mel_filter_coefs[25][104] = 16'h0000;
	mel_filter_coefs[25][105] = 16'h0000;
	mel_filter_coefs[25][106] = 16'h0000;
	mel_filter_coefs[25][107] = 16'h0000;
	mel_filter_coefs[25][108] = 16'h0000;
	mel_filter_coefs[25][109] = 16'h0000;
	mel_filter_coefs[25][110] = 16'h0000;
	mel_filter_coefs[25][111] = 16'h0000;
	mel_filter_coefs[25][112] = 16'h0000;
	mel_filter_coefs[25][113] = 16'h0000;
	mel_filter_coefs[25][114] = 16'h0000;
	mel_filter_coefs[25][115] = 16'h0000;
	mel_filter_coefs[25][116] = 16'h0000;
	mel_filter_coefs[25][117] = 16'h0000;
	mel_filter_coefs[25][118] = 16'h0000;
	mel_filter_coefs[25][119] = 16'h0000;
	mel_filter_coefs[25][120] = 16'h0000;
	mel_filter_coefs[25][121] = 16'h0000;
	mel_filter_coefs[25][122] = 16'h0000;
	mel_filter_coefs[25][123] = 16'h0000;
	mel_filter_coefs[25][124] = 16'h0000;
	mel_filter_coefs[25][125] = 16'h0000;
	mel_filter_coefs[25][126] = 16'h0000;
	mel_filter_coefs[25][127] = 16'h0000;
	mel_filter_coefs[25][128] = 16'h0000;
	mel_filter_coefs[25][129] = 16'h0000;
	mel_filter_coefs[25][130] = 16'h0000;
	mel_filter_coefs[25][131] = 16'h0000;
	mel_filter_coefs[25][132] = 16'h0000;
	mel_filter_coefs[25][133] = 16'h0000;
	mel_filter_coefs[25][134] = 16'h0000;
	mel_filter_coefs[25][135] = 16'h0000;
	mel_filter_coefs[25][136] = 16'h0000;
	mel_filter_coefs[25][137] = 16'h0000;
	mel_filter_coefs[25][138] = 16'h0000;
	mel_filter_coefs[25][139] = 16'h0000;
	mel_filter_coefs[25][140] = 16'h0000;
	mel_filter_coefs[25][141] = 16'h0000;
	mel_filter_coefs[25][142] = 16'h0000;
	mel_filter_coefs[25][143] = 16'h0000;
	mel_filter_coefs[25][144] = 16'h0000;
	mel_filter_coefs[25][145] = 16'h0000;
	mel_filter_coefs[25][146] = 16'h0000;
	mel_filter_coefs[25][147] = 16'h0000;
	mel_filter_coefs[25][148] = 16'h0000;
	mel_filter_coefs[25][149] = 16'h0000;
	mel_filter_coefs[25][150] = 16'h0000;
	mel_filter_coefs[25][151] = 16'h0000;
	mel_filter_coefs[25][152] = 16'h0000;
	mel_filter_coefs[25][153] = 16'h0000;
	mel_filter_coefs[25][154] = 16'h0000;
	mel_filter_coefs[25][155] = 16'h0000;
	mel_filter_coefs[25][156] = 16'h0000;
	mel_filter_coefs[25][157] = 16'h0000;
	mel_filter_coefs[25][158] = 16'h0000;
	mel_filter_coefs[25][159] = 16'h0000;
	mel_filter_coefs[25][160] = 16'h0000;
	mel_filter_coefs[25][161] = 16'h0000;
	mel_filter_coefs[25][162] = 16'h0000;
	mel_filter_coefs[25][163] = 16'h0000;
	mel_filter_coefs[25][164] = 16'h0000;
	mel_filter_coefs[25][165] = 16'h0000;
	mel_filter_coefs[25][166] = 16'h0000;
	mel_filter_coefs[25][167] = 16'h0000;
	mel_filter_coefs[25][168] = 16'h0000;
	mel_filter_coefs[25][169] = 16'h0000;
	mel_filter_coefs[25][170] = 16'h0000;
	mel_filter_coefs[25][171] = 16'h0000;
	mel_filter_coefs[25][172] = 16'h0000;
	mel_filter_coefs[25][173] = 16'h0000;
	mel_filter_coefs[25][174] = 16'h0000;
	mel_filter_coefs[25][175] = 16'h0000;
	mel_filter_coefs[25][176] = 16'h0000;
	mel_filter_coefs[25][177] = 16'h0000;
	mel_filter_coefs[25][178] = 16'h0000;
	mel_filter_coefs[25][179] = 16'h0000;
	mel_filter_coefs[25][180] = 16'h0000;
	mel_filter_coefs[25][181] = 16'h0000;
	mel_filter_coefs[25][182] = 16'h0000;
	mel_filter_coefs[25][183] = 16'h0000;
	mel_filter_coefs[25][184] = 16'h0000;
	mel_filter_coefs[25][185] = 16'h0000;
	mel_filter_coefs[25][186] = 16'h0000;
	mel_filter_coefs[25][187] = 16'h0000;
	mel_filter_coefs[25][188] = 16'h0000;
	mel_filter_coefs[25][189] = 16'h0000;
	mel_filter_coefs[25][190] = 16'h0000;
	mel_filter_coefs[25][191] = 16'h0000;
	mel_filter_coefs[25][192] = 16'h0000;
	mel_filter_coefs[25][193] = 16'h0000;
	mel_filter_coefs[25][194] = 16'h0000;
	mel_filter_coefs[25][195] = 16'h0000;
	mel_filter_coefs[25][196] = 16'h0000;
	mel_filter_coefs[25][197] = 16'h0000;
	mel_filter_coefs[25][198] = 16'h0000;
	mel_filter_coefs[25][199] = 16'h0000;
	mel_filter_coefs[25][200] = 16'h0000;
	mel_filter_coefs[25][201] = 16'h0000;
	mel_filter_coefs[25][202] = 16'h0000;
	mel_filter_coefs[25][203] = 16'h0000;
	mel_filter_coefs[25][204] = 16'h0000;
	mel_filter_coefs[25][205] = 16'h0000;
	mel_filter_coefs[25][206] = 16'h0000;
	mel_filter_coefs[25][207] = 16'h0000;
	mel_filter_coefs[25][208] = 16'h0000;
	mel_filter_coefs[25][209] = 16'h0000;
	mel_filter_coefs[25][210] = 16'h0000;
	mel_filter_coefs[25][211] = 16'h0000;
	mel_filter_coefs[25][212] = 16'h0000;
	mel_filter_coefs[25][213] = 16'h0000;
	mel_filter_coefs[25][214] = 16'h0000;
	mel_filter_coefs[25][215] = 16'h0000;
	mel_filter_coefs[25][216] = 16'h0000;
	mel_filter_coefs[25][217] = 16'h0000;
	mel_filter_coefs[25][218] = 16'h0000;
	mel_filter_coefs[25][219] = 16'h0000;
	mel_filter_coefs[25][220] = 16'h0000;
	mel_filter_coefs[25][221] = 16'h0000;
	mel_filter_coefs[25][222] = 16'h0000;
	mel_filter_coefs[25][223] = 16'h0000;
	mel_filter_coefs[25][224] = 16'h0000;
	mel_filter_coefs[25][225] = 16'h0000;
	mel_filter_coefs[25][226] = 16'h0000;
	mel_filter_coefs[25][227] = 16'h0000;
	mel_filter_coefs[25][228] = 16'h0000;
	mel_filter_coefs[25][229] = 16'h0000;
	mel_filter_coefs[25][230] = 16'h0000;
	mel_filter_coefs[25][231] = 16'h0000;
	mel_filter_coefs[25][232] = 16'h0000;
	mel_filter_coefs[25][233] = 16'h0000;
	mel_filter_coefs[25][234] = 16'h0000;
	mel_filter_coefs[25][235] = 16'h0000;
	mel_filter_coefs[25][236] = 16'h0000;
	mel_filter_coefs[25][237] = 16'h0000;
	mel_filter_coefs[25][238] = 16'h0000;
	mel_filter_coefs[25][239] = 16'h0000;
	mel_filter_coefs[25][240] = 16'h0000;
	mel_filter_coefs[25][241] = 16'h0000;
	mel_filter_coefs[25][242] = 16'h0000;
	mel_filter_coefs[25][243] = 16'h0000;
	mel_filter_coefs[25][244] = 16'h0000;
	mel_filter_coefs[25][245] = 16'h0000;
	mel_filter_coefs[25][246] = 16'h0000;
	mel_filter_coefs[25][247] = 16'h0000;
	mel_filter_coefs[25][248] = 16'h0000;
	mel_filter_coefs[25][249] = 16'h0000;
	mel_filter_coefs[25][250] = 16'h0000;
	mel_filter_coefs[25][251] = 16'h0000;
	mel_filter_coefs[25][252] = 16'h0000;
	mel_filter_coefs[25][253] = 16'h0000;
	mel_filter_coefs[25][254] = 16'h0000;
	mel_filter_coefs[25][255] = 16'h0000;
	mel_filter_coefs[26][0] = 16'h0000;
	mel_filter_coefs[26][1] = 16'h0000;
	mel_filter_coefs[26][2] = 16'h0000;
	mel_filter_coefs[26][3] = 16'h0000;
	mel_filter_coefs[26][4] = 16'h0000;
	mel_filter_coefs[26][5] = 16'h0000;
	mel_filter_coefs[26][6] = 16'h0000;
	mel_filter_coefs[26][7] = 16'h0000;
	mel_filter_coefs[26][8] = 16'h0000;
	mel_filter_coefs[26][9] = 16'h0000;
	mel_filter_coefs[26][10] = 16'h0000;
	mel_filter_coefs[26][11] = 16'h0000;
	mel_filter_coefs[26][12] = 16'h0000;
	mel_filter_coefs[26][13] = 16'h0000;
	mel_filter_coefs[26][14] = 16'h0000;
	mel_filter_coefs[26][15] = 16'h0000;
	mel_filter_coefs[26][16] = 16'h0000;
	mel_filter_coefs[26][17] = 16'h0000;
	mel_filter_coefs[26][18] = 16'h0000;
	mel_filter_coefs[26][19] = 16'h0000;
	mel_filter_coefs[26][20] = 16'h0000;
	mel_filter_coefs[26][21] = 16'h0000;
	mel_filter_coefs[26][22] = 16'h0000;
	mel_filter_coefs[26][23] = 16'h0000;
	mel_filter_coefs[26][24] = 16'h0000;
	mel_filter_coefs[26][25] = 16'h0000;
	mel_filter_coefs[26][26] = 16'h0000;
	mel_filter_coefs[26][27] = 16'h0000;
	mel_filter_coefs[26][28] = 16'h0000;
	mel_filter_coefs[26][29] = 16'h0000;
	mel_filter_coefs[26][30] = 16'h0000;
	mel_filter_coefs[26][31] = 16'h0000;
	mel_filter_coefs[26][32] = 16'h0000;
	mel_filter_coefs[26][33] = 16'h0000;
	mel_filter_coefs[26][34] = 16'h0000;
	mel_filter_coefs[26][35] = 16'h0000;
	mel_filter_coefs[26][36] = 16'h0000;
	mel_filter_coefs[26][37] = 16'h0000;
	mel_filter_coefs[26][38] = 16'h0000;
	mel_filter_coefs[26][39] = 16'h0000;
	mel_filter_coefs[26][40] = 16'h0000;
	mel_filter_coefs[26][41] = 16'h0000;
	mel_filter_coefs[26][42] = 16'h0000;
	mel_filter_coefs[26][43] = 16'h0000;
	mel_filter_coefs[26][44] = 16'h0000;
	mel_filter_coefs[26][45] = 16'h0000;
	mel_filter_coefs[26][46] = 16'h0000;
	mel_filter_coefs[26][47] = 16'h0000;
	mel_filter_coefs[26][48] = 16'h0000;
	mel_filter_coefs[26][49] = 16'h0000;
	mel_filter_coefs[26][50] = 16'h0000;
	mel_filter_coefs[26][51] = 16'h0000;
	mel_filter_coefs[26][52] = 16'h0000;
	mel_filter_coefs[26][53] = 16'h0000;
	mel_filter_coefs[26][54] = 16'h0000;
	mel_filter_coefs[26][55] = 16'h0000;
	mel_filter_coefs[26][56] = 16'h0000;
	mel_filter_coefs[26][57] = 16'h0000;
	mel_filter_coefs[26][58] = 16'h0000;
	mel_filter_coefs[26][59] = 16'h0000;
	mel_filter_coefs[26][60] = 16'h0000;
	mel_filter_coefs[26][61] = 16'h0000;
	mel_filter_coefs[26][62] = 16'h0000;
	mel_filter_coefs[26][63] = 16'h0000;
	mel_filter_coefs[26][64] = 16'h0000;
	mel_filter_coefs[26][65] = 16'h0000;
	mel_filter_coefs[26][66] = 16'h0000;
	mel_filter_coefs[26][67] = 16'h0000;
	mel_filter_coefs[26][68] = 16'h0000;
	mel_filter_coefs[26][69] = 16'h0000;
	mel_filter_coefs[26][70] = 16'h0000;
	mel_filter_coefs[26][71] = 16'h0000;
	mel_filter_coefs[26][72] = 16'h0000;
	mel_filter_coefs[26][73] = 16'h0000;
	mel_filter_coefs[26][74] = 16'h0000;
	mel_filter_coefs[26][75] = 16'h0000;
	mel_filter_coefs[26][76] = 16'h0000;
	mel_filter_coefs[26][77] = 16'h0000;
	mel_filter_coefs[26][78] = 16'h0000;
	mel_filter_coefs[26][79] = 16'h0000;
	mel_filter_coefs[26][80] = 16'h0000;
	mel_filter_coefs[26][81] = 16'h0000;
	mel_filter_coefs[26][82] = 16'h0000;
	mel_filter_coefs[26][83] = 16'h0000;
	mel_filter_coefs[26][84] = 16'h0000;
	mel_filter_coefs[26][85] = 16'h0000;
	mel_filter_coefs[26][86] = 16'h0000;
	mel_filter_coefs[26][87] = 16'h0000;
	mel_filter_coefs[26][88] = 16'h003F;
	mel_filter_coefs[26][89] = 16'h128E;
	mel_filter_coefs[26][90] = 16'h24DC;
	mel_filter_coefs[26][91] = 16'h372B;
	mel_filter_coefs[26][92] = 16'h4979;
	mel_filter_coefs[26][93] = 16'h5BC8;
	mel_filter_coefs[26][94] = 16'h6E16;
	mel_filter_coefs[26][95] = 16'h7FA1;
	mel_filter_coefs[26][96] = 16'h6E6A;
	mel_filter_coefs[26][97] = 16'h5D33;
	mel_filter_coefs[26][98] = 16'h4BFC;
	mel_filter_coefs[26][99] = 16'h3AC5;
	mel_filter_coefs[26][100] = 16'h298E;
	mel_filter_coefs[26][101] = 16'h1857;
	mel_filter_coefs[26][102] = 16'h071F;
	mel_filter_coefs[26][103] = 16'h0000;
	mel_filter_coefs[26][104] = 16'h0000;
	mel_filter_coefs[26][105] = 16'h0000;
	mel_filter_coefs[26][106] = 16'h0000;
	mel_filter_coefs[26][107] = 16'h0000;
	mel_filter_coefs[26][108] = 16'h0000;
	mel_filter_coefs[26][109] = 16'h0000;
	mel_filter_coefs[26][110] = 16'h0000;
	mel_filter_coefs[26][111] = 16'h0000;
	mel_filter_coefs[26][112] = 16'h0000;
	mel_filter_coefs[26][113] = 16'h0000;
	mel_filter_coefs[26][114] = 16'h0000;
	mel_filter_coefs[26][115] = 16'h0000;
	mel_filter_coefs[26][116] = 16'h0000;
	mel_filter_coefs[26][117] = 16'h0000;
	mel_filter_coefs[26][118] = 16'h0000;
	mel_filter_coefs[26][119] = 16'h0000;
	mel_filter_coefs[26][120] = 16'h0000;
	mel_filter_coefs[26][121] = 16'h0000;
	mel_filter_coefs[26][122] = 16'h0000;
	mel_filter_coefs[26][123] = 16'h0000;
	mel_filter_coefs[26][124] = 16'h0000;
	mel_filter_coefs[26][125] = 16'h0000;
	mel_filter_coefs[26][126] = 16'h0000;
	mel_filter_coefs[26][127] = 16'h0000;
	mel_filter_coefs[26][128] = 16'h0000;
	mel_filter_coefs[26][129] = 16'h0000;
	mel_filter_coefs[26][130] = 16'h0000;
	mel_filter_coefs[26][131] = 16'h0000;
	mel_filter_coefs[26][132] = 16'h0000;
	mel_filter_coefs[26][133] = 16'h0000;
	mel_filter_coefs[26][134] = 16'h0000;
	mel_filter_coefs[26][135] = 16'h0000;
	mel_filter_coefs[26][136] = 16'h0000;
	mel_filter_coefs[26][137] = 16'h0000;
	mel_filter_coefs[26][138] = 16'h0000;
	mel_filter_coefs[26][139] = 16'h0000;
	mel_filter_coefs[26][140] = 16'h0000;
	mel_filter_coefs[26][141] = 16'h0000;
	mel_filter_coefs[26][142] = 16'h0000;
	mel_filter_coefs[26][143] = 16'h0000;
	mel_filter_coefs[26][144] = 16'h0000;
	mel_filter_coefs[26][145] = 16'h0000;
	mel_filter_coefs[26][146] = 16'h0000;
	mel_filter_coefs[26][147] = 16'h0000;
	mel_filter_coefs[26][148] = 16'h0000;
	mel_filter_coefs[26][149] = 16'h0000;
	mel_filter_coefs[26][150] = 16'h0000;
	mel_filter_coefs[26][151] = 16'h0000;
	mel_filter_coefs[26][152] = 16'h0000;
	mel_filter_coefs[26][153] = 16'h0000;
	mel_filter_coefs[26][154] = 16'h0000;
	mel_filter_coefs[26][155] = 16'h0000;
	mel_filter_coefs[26][156] = 16'h0000;
	mel_filter_coefs[26][157] = 16'h0000;
	mel_filter_coefs[26][158] = 16'h0000;
	mel_filter_coefs[26][159] = 16'h0000;
	mel_filter_coefs[26][160] = 16'h0000;
	mel_filter_coefs[26][161] = 16'h0000;
	mel_filter_coefs[26][162] = 16'h0000;
	mel_filter_coefs[26][163] = 16'h0000;
	mel_filter_coefs[26][164] = 16'h0000;
	mel_filter_coefs[26][165] = 16'h0000;
	mel_filter_coefs[26][166] = 16'h0000;
	mel_filter_coefs[26][167] = 16'h0000;
	mel_filter_coefs[26][168] = 16'h0000;
	mel_filter_coefs[26][169] = 16'h0000;
	mel_filter_coefs[26][170] = 16'h0000;
	mel_filter_coefs[26][171] = 16'h0000;
	mel_filter_coefs[26][172] = 16'h0000;
	mel_filter_coefs[26][173] = 16'h0000;
	mel_filter_coefs[26][174] = 16'h0000;
	mel_filter_coefs[26][175] = 16'h0000;
	mel_filter_coefs[26][176] = 16'h0000;
	mel_filter_coefs[26][177] = 16'h0000;
	mel_filter_coefs[26][178] = 16'h0000;
	mel_filter_coefs[26][179] = 16'h0000;
	mel_filter_coefs[26][180] = 16'h0000;
	mel_filter_coefs[26][181] = 16'h0000;
	mel_filter_coefs[26][182] = 16'h0000;
	mel_filter_coefs[26][183] = 16'h0000;
	mel_filter_coefs[26][184] = 16'h0000;
	mel_filter_coefs[26][185] = 16'h0000;
	mel_filter_coefs[26][186] = 16'h0000;
	mel_filter_coefs[26][187] = 16'h0000;
	mel_filter_coefs[26][188] = 16'h0000;
	mel_filter_coefs[26][189] = 16'h0000;
	mel_filter_coefs[26][190] = 16'h0000;
	mel_filter_coefs[26][191] = 16'h0000;
	mel_filter_coefs[26][192] = 16'h0000;
	mel_filter_coefs[26][193] = 16'h0000;
	mel_filter_coefs[26][194] = 16'h0000;
	mel_filter_coefs[26][195] = 16'h0000;
	mel_filter_coefs[26][196] = 16'h0000;
	mel_filter_coefs[26][197] = 16'h0000;
	mel_filter_coefs[26][198] = 16'h0000;
	mel_filter_coefs[26][199] = 16'h0000;
	mel_filter_coefs[26][200] = 16'h0000;
	mel_filter_coefs[26][201] = 16'h0000;
	mel_filter_coefs[26][202] = 16'h0000;
	mel_filter_coefs[26][203] = 16'h0000;
	mel_filter_coefs[26][204] = 16'h0000;
	mel_filter_coefs[26][205] = 16'h0000;
	mel_filter_coefs[26][206] = 16'h0000;
	mel_filter_coefs[26][207] = 16'h0000;
	mel_filter_coefs[26][208] = 16'h0000;
	mel_filter_coefs[26][209] = 16'h0000;
	mel_filter_coefs[26][210] = 16'h0000;
	mel_filter_coefs[26][211] = 16'h0000;
	mel_filter_coefs[26][212] = 16'h0000;
	mel_filter_coefs[26][213] = 16'h0000;
	mel_filter_coefs[26][214] = 16'h0000;
	mel_filter_coefs[26][215] = 16'h0000;
	mel_filter_coefs[26][216] = 16'h0000;
	mel_filter_coefs[26][217] = 16'h0000;
	mel_filter_coefs[26][218] = 16'h0000;
	mel_filter_coefs[26][219] = 16'h0000;
	mel_filter_coefs[26][220] = 16'h0000;
	mel_filter_coefs[26][221] = 16'h0000;
	mel_filter_coefs[26][222] = 16'h0000;
	mel_filter_coefs[26][223] = 16'h0000;
	mel_filter_coefs[26][224] = 16'h0000;
	mel_filter_coefs[26][225] = 16'h0000;
	mel_filter_coefs[26][226] = 16'h0000;
	mel_filter_coefs[26][227] = 16'h0000;
	mel_filter_coefs[26][228] = 16'h0000;
	mel_filter_coefs[26][229] = 16'h0000;
	mel_filter_coefs[26][230] = 16'h0000;
	mel_filter_coefs[26][231] = 16'h0000;
	mel_filter_coefs[26][232] = 16'h0000;
	mel_filter_coefs[26][233] = 16'h0000;
	mel_filter_coefs[26][234] = 16'h0000;
	mel_filter_coefs[26][235] = 16'h0000;
	mel_filter_coefs[26][236] = 16'h0000;
	mel_filter_coefs[26][237] = 16'h0000;
	mel_filter_coefs[26][238] = 16'h0000;
	mel_filter_coefs[26][239] = 16'h0000;
	mel_filter_coefs[26][240] = 16'h0000;
	mel_filter_coefs[26][241] = 16'h0000;
	mel_filter_coefs[26][242] = 16'h0000;
	mel_filter_coefs[26][243] = 16'h0000;
	mel_filter_coefs[26][244] = 16'h0000;
	mel_filter_coefs[26][245] = 16'h0000;
	mel_filter_coefs[26][246] = 16'h0000;
	mel_filter_coefs[26][247] = 16'h0000;
	mel_filter_coefs[26][248] = 16'h0000;
	mel_filter_coefs[26][249] = 16'h0000;
	mel_filter_coefs[26][250] = 16'h0000;
	mel_filter_coefs[26][251] = 16'h0000;
	mel_filter_coefs[26][252] = 16'h0000;
	mel_filter_coefs[26][253] = 16'h0000;
	mel_filter_coefs[26][254] = 16'h0000;
	mel_filter_coefs[26][255] = 16'h0000;
	mel_filter_coefs[27][0] = 16'h0000;
	mel_filter_coefs[27][1] = 16'h0000;
	mel_filter_coefs[27][2] = 16'h0000;
	mel_filter_coefs[27][3] = 16'h0000;
	mel_filter_coefs[27][4] = 16'h0000;
	mel_filter_coefs[27][5] = 16'h0000;
	mel_filter_coefs[27][6] = 16'h0000;
	mel_filter_coefs[27][7] = 16'h0000;
	mel_filter_coefs[27][8] = 16'h0000;
	mel_filter_coefs[27][9] = 16'h0000;
	mel_filter_coefs[27][10] = 16'h0000;
	mel_filter_coefs[27][11] = 16'h0000;
	mel_filter_coefs[27][12] = 16'h0000;
	mel_filter_coefs[27][13] = 16'h0000;
	mel_filter_coefs[27][14] = 16'h0000;
	mel_filter_coefs[27][15] = 16'h0000;
	mel_filter_coefs[27][16] = 16'h0000;
	mel_filter_coefs[27][17] = 16'h0000;
	mel_filter_coefs[27][18] = 16'h0000;
	mel_filter_coefs[27][19] = 16'h0000;
	mel_filter_coefs[27][20] = 16'h0000;
	mel_filter_coefs[27][21] = 16'h0000;
	mel_filter_coefs[27][22] = 16'h0000;
	mel_filter_coefs[27][23] = 16'h0000;
	mel_filter_coefs[27][24] = 16'h0000;
	mel_filter_coefs[27][25] = 16'h0000;
	mel_filter_coefs[27][26] = 16'h0000;
	mel_filter_coefs[27][27] = 16'h0000;
	mel_filter_coefs[27][28] = 16'h0000;
	mel_filter_coefs[27][29] = 16'h0000;
	mel_filter_coefs[27][30] = 16'h0000;
	mel_filter_coefs[27][31] = 16'h0000;
	mel_filter_coefs[27][32] = 16'h0000;
	mel_filter_coefs[27][33] = 16'h0000;
	mel_filter_coefs[27][34] = 16'h0000;
	mel_filter_coefs[27][35] = 16'h0000;
	mel_filter_coefs[27][36] = 16'h0000;
	mel_filter_coefs[27][37] = 16'h0000;
	mel_filter_coefs[27][38] = 16'h0000;
	mel_filter_coefs[27][39] = 16'h0000;
	mel_filter_coefs[27][40] = 16'h0000;
	mel_filter_coefs[27][41] = 16'h0000;
	mel_filter_coefs[27][42] = 16'h0000;
	mel_filter_coefs[27][43] = 16'h0000;
	mel_filter_coefs[27][44] = 16'h0000;
	mel_filter_coefs[27][45] = 16'h0000;
	mel_filter_coefs[27][46] = 16'h0000;
	mel_filter_coefs[27][47] = 16'h0000;
	mel_filter_coefs[27][48] = 16'h0000;
	mel_filter_coefs[27][49] = 16'h0000;
	mel_filter_coefs[27][50] = 16'h0000;
	mel_filter_coefs[27][51] = 16'h0000;
	mel_filter_coefs[27][52] = 16'h0000;
	mel_filter_coefs[27][53] = 16'h0000;
	mel_filter_coefs[27][54] = 16'h0000;
	mel_filter_coefs[27][55] = 16'h0000;
	mel_filter_coefs[27][56] = 16'h0000;
	mel_filter_coefs[27][57] = 16'h0000;
	mel_filter_coefs[27][58] = 16'h0000;
	mel_filter_coefs[27][59] = 16'h0000;
	mel_filter_coefs[27][60] = 16'h0000;
	mel_filter_coefs[27][61] = 16'h0000;
	mel_filter_coefs[27][62] = 16'h0000;
	mel_filter_coefs[27][63] = 16'h0000;
	mel_filter_coefs[27][64] = 16'h0000;
	mel_filter_coefs[27][65] = 16'h0000;
	mel_filter_coefs[27][66] = 16'h0000;
	mel_filter_coefs[27][67] = 16'h0000;
	mel_filter_coefs[27][68] = 16'h0000;
	mel_filter_coefs[27][69] = 16'h0000;
	mel_filter_coefs[27][70] = 16'h0000;
	mel_filter_coefs[27][71] = 16'h0000;
	mel_filter_coefs[27][72] = 16'h0000;
	mel_filter_coefs[27][73] = 16'h0000;
	mel_filter_coefs[27][74] = 16'h0000;
	mel_filter_coefs[27][75] = 16'h0000;
	mel_filter_coefs[27][76] = 16'h0000;
	mel_filter_coefs[27][77] = 16'h0000;
	mel_filter_coefs[27][78] = 16'h0000;
	mel_filter_coefs[27][79] = 16'h0000;
	mel_filter_coefs[27][80] = 16'h0000;
	mel_filter_coefs[27][81] = 16'h0000;
	mel_filter_coefs[27][82] = 16'h0000;
	mel_filter_coefs[27][83] = 16'h0000;
	mel_filter_coefs[27][84] = 16'h0000;
	mel_filter_coefs[27][85] = 16'h0000;
	mel_filter_coefs[27][86] = 16'h0000;
	mel_filter_coefs[27][87] = 16'h0000;
	mel_filter_coefs[27][88] = 16'h0000;
	mel_filter_coefs[27][89] = 16'h0000;
	mel_filter_coefs[27][90] = 16'h0000;
	mel_filter_coefs[27][91] = 16'h0000;
	mel_filter_coefs[27][92] = 16'h0000;
	mel_filter_coefs[27][93] = 16'h0000;
	mel_filter_coefs[27][94] = 16'h0000;
	mel_filter_coefs[27][95] = 16'h005F;
	mel_filter_coefs[27][96] = 16'h1196;
	mel_filter_coefs[27][97] = 16'h22CD;
	mel_filter_coefs[27][98] = 16'h3404;
	mel_filter_coefs[27][99] = 16'h453B;
	mel_filter_coefs[27][100] = 16'h5672;
	mel_filter_coefs[27][101] = 16'h67A9;
	mel_filter_coefs[27][102] = 16'h78E1;
	mel_filter_coefs[27][103] = 16'h7682;
	mel_filter_coefs[27][104] = 16'h6652;
	mel_filter_coefs[27][105] = 16'h5622;
	mel_filter_coefs[27][106] = 16'h45F1;
	mel_filter_coefs[27][107] = 16'h35C1;
	mel_filter_coefs[27][108] = 16'h2590;
	mel_filter_coefs[27][109] = 16'h1560;
	mel_filter_coefs[27][110] = 16'h0530;
	mel_filter_coefs[27][111] = 16'h0000;
	mel_filter_coefs[27][112] = 16'h0000;
	mel_filter_coefs[27][113] = 16'h0000;
	mel_filter_coefs[27][114] = 16'h0000;
	mel_filter_coefs[27][115] = 16'h0000;
	mel_filter_coefs[27][116] = 16'h0000;
	mel_filter_coefs[27][117] = 16'h0000;
	mel_filter_coefs[27][118] = 16'h0000;
	mel_filter_coefs[27][119] = 16'h0000;
	mel_filter_coefs[27][120] = 16'h0000;
	mel_filter_coefs[27][121] = 16'h0000;
	mel_filter_coefs[27][122] = 16'h0000;
	mel_filter_coefs[27][123] = 16'h0000;
	mel_filter_coefs[27][124] = 16'h0000;
	mel_filter_coefs[27][125] = 16'h0000;
	mel_filter_coefs[27][126] = 16'h0000;
	mel_filter_coefs[27][127] = 16'h0000;
	mel_filter_coefs[27][128] = 16'h0000;
	mel_filter_coefs[27][129] = 16'h0000;
	mel_filter_coefs[27][130] = 16'h0000;
	mel_filter_coefs[27][131] = 16'h0000;
	mel_filter_coefs[27][132] = 16'h0000;
	mel_filter_coefs[27][133] = 16'h0000;
	mel_filter_coefs[27][134] = 16'h0000;
	mel_filter_coefs[27][135] = 16'h0000;
	mel_filter_coefs[27][136] = 16'h0000;
	mel_filter_coefs[27][137] = 16'h0000;
	mel_filter_coefs[27][138] = 16'h0000;
	mel_filter_coefs[27][139] = 16'h0000;
	mel_filter_coefs[27][140] = 16'h0000;
	mel_filter_coefs[27][141] = 16'h0000;
	mel_filter_coefs[27][142] = 16'h0000;
	mel_filter_coefs[27][143] = 16'h0000;
	mel_filter_coefs[27][144] = 16'h0000;
	mel_filter_coefs[27][145] = 16'h0000;
	mel_filter_coefs[27][146] = 16'h0000;
	mel_filter_coefs[27][147] = 16'h0000;
	mel_filter_coefs[27][148] = 16'h0000;
	mel_filter_coefs[27][149] = 16'h0000;
	mel_filter_coefs[27][150] = 16'h0000;
	mel_filter_coefs[27][151] = 16'h0000;
	mel_filter_coefs[27][152] = 16'h0000;
	mel_filter_coefs[27][153] = 16'h0000;
	mel_filter_coefs[27][154] = 16'h0000;
	mel_filter_coefs[27][155] = 16'h0000;
	mel_filter_coefs[27][156] = 16'h0000;
	mel_filter_coefs[27][157] = 16'h0000;
	mel_filter_coefs[27][158] = 16'h0000;
	mel_filter_coefs[27][159] = 16'h0000;
	mel_filter_coefs[27][160] = 16'h0000;
	mel_filter_coefs[27][161] = 16'h0000;
	mel_filter_coefs[27][162] = 16'h0000;
	mel_filter_coefs[27][163] = 16'h0000;
	mel_filter_coefs[27][164] = 16'h0000;
	mel_filter_coefs[27][165] = 16'h0000;
	mel_filter_coefs[27][166] = 16'h0000;
	mel_filter_coefs[27][167] = 16'h0000;
	mel_filter_coefs[27][168] = 16'h0000;
	mel_filter_coefs[27][169] = 16'h0000;
	mel_filter_coefs[27][170] = 16'h0000;
	mel_filter_coefs[27][171] = 16'h0000;
	mel_filter_coefs[27][172] = 16'h0000;
	mel_filter_coefs[27][173] = 16'h0000;
	mel_filter_coefs[27][174] = 16'h0000;
	mel_filter_coefs[27][175] = 16'h0000;
	mel_filter_coefs[27][176] = 16'h0000;
	mel_filter_coefs[27][177] = 16'h0000;
	mel_filter_coefs[27][178] = 16'h0000;
	mel_filter_coefs[27][179] = 16'h0000;
	mel_filter_coefs[27][180] = 16'h0000;
	mel_filter_coefs[27][181] = 16'h0000;
	mel_filter_coefs[27][182] = 16'h0000;
	mel_filter_coefs[27][183] = 16'h0000;
	mel_filter_coefs[27][184] = 16'h0000;
	mel_filter_coefs[27][185] = 16'h0000;
	mel_filter_coefs[27][186] = 16'h0000;
	mel_filter_coefs[27][187] = 16'h0000;
	mel_filter_coefs[27][188] = 16'h0000;
	mel_filter_coefs[27][189] = 16'h0000;
	mel_filter_coefs[27][190] = 16'h0000;
	mel_filter_coefs[27][191] = 16'h0000;
	mel_filter_coefs[27][192] = 16'h0000;
	mel_filter_coefs[27][193] = 16'h0000;
	mel_filter_coefs[27][194] = 16'h0000;
	mel_filter_coefs[27][195] = 16'h0000;
	mel_filter_coefs[27][196] = 16'h0000;
	mel_filter_coefs[27][197] = 16'h0000;
	mel_filter_coefs[27][198] = 16'h0000;
	mel_filter_coefs[27][199] = 16'h0000;
	mel_filter_coefs[27][200] = 16'h0000;
	mel_filter_coefs[27][201] = 16'h0000;
	mel_filter_coefs[27][202] = 16'h0000;
	mel_filter_coefs[27][203] = 16'h0000;
	mel_filter_coefs[27][204] = 16'h0000;
	mel_filter_coefs[27][205] = 16'h0000;
	mel_filter_coefs[27][206] = 16'h0000;
	mel_filter_coefs[27][207] = 16'h0000;
	mel_filter_coefs[27][208] = 16'h0000;
	mel_filter_coefs[27][209] = 16'h0000;
	mel_filter_coefs[27][210] = 16'h0000;
	mel_filter_coefs[27][211] = 16'h0000;
	mel_filter_coefs[27][212] = 16'h0000;
	mel_filter_coefs[27][213] = 16'h0000;
	mel_filter_coefs[27][214] = 16'h0000;
	mel_filter_coefs[27][215] = 16'h0000;
	mel_filter_coefs[27][216] = 16'h0000;
	mel_filter_coefs[27][217] = 16'h0000;
	mel_filter_coefs[27][218] = 16'h0000;
	mel_filter_coefs[27][219] = 16'h0000;
	mel_filter_coefs[27][220] = 16'h0000;
	mel_filter_coefs[27][221] = 16'h0000;
	mel_filter_coefs[27][222] = 16'h0000;
	mel_filter_coefs[27][223] = 16'h0000;
	mel_filter_coefs[27][224] = 16'h0000;
	mel_filter_coefs[27][225] = 16'h0000;
	mel_filter_coefs[27][226] = 16'h0000;
	mel_filter_coefs[27][227] = 16'h0000;
	mel_filter_coefs[27][228] = 16'h0000;
	mel_filter_coefs[27][229] = 16'h0000;
	mel_filter_coefs[27][230] = 16'h0000;
	mel_filter_coefs[27][231] = 16'h0000;
	mel_filter_coefs[27][232] = 16'h0000;
	mel_filter_coefs[27][233] = 16'h0000;
	mel_filter_coefs[27][234] = 16'h0000;
	mel_filter_coefs[27][235] = 16'h0000;
	mel_filter_coefs[27][236] = 16'h0000;
	mel_filter_coefs[27][237] = 16'h0000;
	mel_filter_coefs[27][238] = 16'h0000;
	mel_filter_coefs[27][239] = 16'h0000;
	mel_filter_coefs[27][240] = 16'h0000;
	mel_filter_coefs[27][241] = 16'h0000;
	mel_filter_coefs[27][242] = 16'h0000;
	mel_filter_coefs[27][243] = 16'h0000;
	mel_filter_coefs[27][244] = 16'h0000;
	mel_filter_coefs[27][245] = 16'h0000;
	mel_filter_coefs[27][246] = 16'h0000;
	mel_filter_coefs[27][247] = 16'h0000;
	mel_filter_coefs[27][248] = 16'h0000;
	mel_filter_coefs[27][249] = 16'h0000;
	mel_filter_coefs[27][250] = 16'h0000;
	mel_filter_coefs[27][251] = 16'h0000;
	mel_filter_coefs[27][252] = 16'h0000;
	mel_filter_coefs[27][253] = 16'h0000;
	mel_filter_coefs[27][254] = 16'h0000;
	mel_filter_coefs[27][255] = 16'h0000;
	mel_filter_coefs[28][0] = 16'h0000;
	mel_filter_coefs[28][1] = 16'h0000;
	mel_filter_coefs[28][2] = 16'h0000;
	mel_filter_coefs[28][3] = 16'h0000;
	mel_filter_coefs[28][4] = 16'h0000;
	mel_filter_coefs[28][5] = 16'h0000;
	mel_filter_coefs[28][6] = 16'h0000;
	mel_filter_coefs[28][7] = 16'h0000;
	mel_filter_coefs[28][8] = 16'h0000;
	mel_filter_coefs[28][9] = 16'h0000;
	mel_filter_coefs[28][10] = 16'h0000;
	mel_filter_coefs[28][11] = 16'h0000;
	mel_filter_coefs[28][12] = 16'h0000;
	mel_filter_coefs[28][13] = 16'h0000;
	mel_filter_coefs[28][14] = 16'h0000;
	mel_filter_coefs[28][15] = 16'h0000;
	mel_filter_coefs[28][16] = 16'h0000;
	mel_filter_coefs[28][17] = 16'h0000;
	mel_filter_coefs[28][18] = 16'h0000;
	mel_filter_coefs[28][19] = 16'h0000;
	mel_filter_coefs[28][20] = 16'h0000;
	mel_filter_coefs[28][21] = 16'h0000;
	mel_filter_coefs[28][22] = 16'h0000;
	mel_filter_coefs[28][23] = 16'h0000;
	mel_filter_coefs[28][24] = 16'h0000;
	mel_filter_coefs[28][25] = 16'h0000;
	mel_filter_coefs[28][26] = 16'h0000;
	mel_filter_coefs[28][27] = 16'h0000;
	mel_filter_coefs[28][28] = 16'h0000;
	mel_filter_coefs[28][29] = 16'h0000;
	mel_filter_coefs[28][30] = 16'h0000;
	mel_filter_coefs[28][31] = 16'h0000;
	mel_filter_coefs[28][32] = 16'h0000;
	mel_filter_coefs[28][33] = 16'h0000;
	mel_filter_coefs[28][34] = 16'h0000;
	mel_filter_coefs[28][35] = 16'h0000;
	mel_filter_coefs[28][36] = 16'h0000;
	mel_filter_coefs[28][37] = 16'h0000;
	mel_filter_coefs[28][38] = 16'h0000;
	mel_filter_coefs[28][39] = 16'h0000;
	mel_filter_coefs[28][40] = 16'h0000;
	mel_filter_coefs[28][41] = 16'h0000;
	mel_filter_coefs[28][42] = 16'h0000;
	mel_filter_coefs[28][43] = 16'h0000;
	mel_filter_coefs[28][44] = 16'h0000;
	mel_filter_coefs[28][45] = 16'h0000;
	mel_filter_coefs[28][46] = 16'h0000;
	mel_filter_coefs[28][47] = 16'h0000;
	mel_filter_coefs[28][48] = 16'h0000;
	mel_filter_coefs[28][49] = 16'h0000;
	mel_filter_coefs[28][50] = 16'h0000;
	mel_filter_coefs[28][51] = 16'h0000;
	mel_filter_coefs[28][52] = 16'h0000;
	mel_filter_coefs[28][53] = 16'h0000;
	mel_filter_coefs[28][54] = 16'h0000;
	mel_filter_coefs[28][55] = 16'h0000;
	mel_filter_coefs[28][56] = 16'h0000;
	mel_filter_coefs[28][57] = 16'h0000;
	mel_filter_coefs[28][58] = 16'h0000;
	mel_filter_coefs[28][59] = 16'h0000;
	mel_filter_coefs[28][60] = 16'h0000;
	mel_filter_coefs[28][61] = 16'h0000;
	mel_filter_coefs[28][62] = 16'h0000;
	mel_filter_coefs[28][63] = 16'h0000;
	mel_filter_coefs[28][64] = 16'h0000;
	mel_filter_coefs[28][65] = 16'h0000;
	mel_filter_coefs[28][66] = 16'h0000;
	mel_filter_coefs[28][67] = 16'h0000;
	mel_filter_coefs[28][68] = 16'h0000;
	mel_filter_coefs[28][69] = 16'h0000;
	mel_filter_coefs[28][70] = 16'h0000;
	mel_filter_coefs[28][71] = 16'h0000;
	mel_filter_coefs[28][72] = 16'h0000;
	mel_filter_coefs[28][73] = 16'h0000;
	mel_filter_coefs[28][74] = 16'h0000;
	mel_filter_coefs[28][75] = 16'h0000;
	mel_filter_coefs[28][76] = 16'h0000;
	mel_filter_coefs[28][77] = 16'h0000;
	mel_filter_coefs[28][78] = 16'h0000;
	mel_filter_coefs[28][79] = 16'h0000;
	mel_filter_coefs[28][80] = 16'h0000;
	mel_filter_coefs[28][81] = 16'h0000;
	mel_filter_coefs[28][82] = 16'h0000;
	mel_filter_coefs[28][83] = 16'h0000;
	mel_filter_coefs[28][84] = 16'h0000;
	mel_filter_coefs[28][85] = 16'h0000;
	mel_filter_coefs[28][86] = 16'h0000;
	mel_filter_coefs[28][87] = 16'h0000;
	mel_filter_coefs[28][88] = 16'h0000;
	mel_filter_coefs[28][89] = 16'h0000;
	mel_filter_coefs[28][90] = 16'h0000;
	mel_filter_coefs[28][91] = 16'h0000;
	mel_filter_coefs[28][92] = 16'h0000;
	mel_filter_coefs[28][93] = 16'h0000;
	mel_filter_coefs[28][94] = 16'h0000;
	mel_filter_coefs[28][95] = 16'h0000;
	mel_filter_coefs[28][96] = 16'h0000;
	mel_filter_coefs[28][97] = 16'h0000;
	mel_filter_coefs[28][98] = 16'h0000;
	mel_filter_coefs[28][99] = 16'h0000;
	mel_filter_coefs[28][100] = 16'h0000;
	mel_filter_coefs[28][101] = 16'h0000;
	mel_filter_coefs[28][102] = 16'h0000;
	mel_filter_coefs[28][103] = 16'h097E;
	mel_filter_coefs[28][104] = 16'h19AE;
	mel_filter_coefs[28][105] = 16'h29DE;
	mel_filter_coefs[28][106] = 16'h3A0F;
	mel_filter_coefs[28][107] = 16'h4A3F;
	mel_filter_coefs[28][108] = 16'h5A70;
	mel_filter_coefs[28][109] = 16'h6AA0;
	mel_filter_coefs[28][110] = 16'h7AD0;
	mel_filter_coefs[28][111] = 16'h75A7;
	mel_filter_coefs[28][112] = 16'h666E;
	mel_filter_coefs[28][113] = 16'h5734;
	mel_filter_coefs[28][114] = 16'h47FB;
	mel_filter_coefs[28][115] = 16'h38C2;
	mel_filter_coefs[28][116] = 16'h2988;
	mel_filter_coefs[28][117] = 16'h1A4F;
	mel_filter_coefs[28][118] = 16'h0B16;
	mel_filter_coefs[28][119] = 16'h0000;
	mel_filter_coefs[28][120] = 16'h0000;
	mel_filter_coefs[28][121] = 16'h0000;
	mel_filter_coefs[28][122] = 16'h0000;
	mel_filter_coefs[28][123] = 16'h0000;
	mel_filter_coefs[28][124] = 16'h0000;
	mel_filter_coefs[28][125] = 16'h0000;
	mel_filter_coefs[28][126] = 16'h0000;
	mel_filter_coefs[28][127] = 16'h0000;
	mel_filter_coefs[28][128] = 16'h0000;
	mel_filter_coefs[28][129] = 16'h0000;
	mel_filter_coefs[28][130] = 16'h0000;
	mel_filter_coefs[28][131] = 16'h0000;
	mel_filter_coefs[28][132] = 16'h0000;
	mel_filter_coefs[28][133] = 16'h0000;
	mel_filter_coefs[28][134] = 16'h0000;
	mel_filter_coefs[28][135] = 16'h0000;
	mel_filter_coefs[28][136] = 16'h0000;
	mel_filter_coefs[28][137] = 16'h0000;
	mel_filter_coefs[28][138] = 16'h0000;
	mel_filter_coefs[28][139] = 16'h0000;
	mel_filter_coefs[28][140] = 16'h0000;
	mel_filter_coefs[28][141] = 16'h0000;
	mel_filter_coefs[28][142] = 16'h0000;
	mel_filter_coefs[28][143] = 16'h0000;
	mel_filter_coefs[28][144] = 16'h0000;
	mel_filter_coefs[28][145] = 16'h0000;
	mel_filter_coefs[28][146] = 16'h0000;
	mel_filter_coefs[28][147] = 16'h0000;
	mel_filter_coefs[28][148] = 16'h0000;
	mel_filter_coefs[28][149] = 16'h0000;
	mel_filter_coefs[28][150] = 16'h0000;
	mel_filter_coefs[28][151] = 16'h0000;
	mel_filter_coefs[28][152] = 16'h0000;
	mel_filter_coefs[28][153] = 16'h0000;
	mel_filter_coefs[28][154] = 16'h0000;
	mel_filter_coefs[28][155] = 16'h0000;
	mel_filter_coefs[28][156] = 16'h0000;
	mel_filter_coefs[28][157] = 16'h0000;
	mel_filter_coefs[28][158] = 16'h0000;
	mel_filter_coefs[28][159] = 16'h0000;
	mel_filter_coefs[28][160] = 16'h0000;
	mel_filter_coefs[28][161] = 16'h0000;
	mel_filter_coefs[28][162] = 16'h0000;
	mel_filter_coefs[28][163] = 16'h0000;
	mel_filter_coefs[28][164] = 16'h0000;
	mel_filter_coefs[28][165] = 16'h0000;
	mel_filter_coefs[28][166] = 16'h0000;
	mel_filter_coefs[28][167] = 16'h0000;
	mel_filter_coefs[28][168] = 16'h0000;
	mel_filter_coefs[28][169] = 16'h0000;
	mel_filter_coefs[28][170] = 16'h0000;
	mel_filter_coefs[28][171] = 16'h0000;
	mel_filter_coefs[28][172] = 16'h0000;
	mel_filter_coefs[28][173] = 16'h0000;
	mel_filter_coefs[28][174] = 16'h0000;
	mel_filter_coefs[28][175] = 16'h0000;
	mel_filter_coefs[28][176] = 16'h0000;
	mel_filter_coefs[28][177] = 16'h0000;
	mel_filter_coefs[28][178] = 16'h0000;
	mel_filter_coefs[28][179] = 16'h0000;
	mel_filter_coefs[28][180] = 16'h0000;
	mel_filter_coefs[28][181] = 16'h0000;
	mel_filter_coefs[28][182] = 16'h0000;
	mel_filter_coefs[28][183] = 16'h0000;
	mel_filter_coefs[28][184] = 16'h0000;
	mel_filter_coefs[28][185] = 16'h0000;
	mel_filter_coefs[28][186] = 16'h0000;
	mel_filter_coefs[28][187] = 16'h0000;
	mel_filter_coefs[28][188] = 16'h0000;
	mel_filter_coefs[28][189] = 16'h0000;
	mel_filter_coefs[28][190] = 16'h0000;
	mel_filter_coefs[28][191] = 16'h0000;
	mel_filter_coefs[28][192] = 16'h0000;
	mel_filter_coefs[28][193] = 16'h0000;
	mel_filter_coefs[28][194] = 16'h0000;
	mel_filter_coefs[28][195] = 16'h0000;
	mel_filter_coefs[28][196] = 16'h0000;
	mel_filter_coefs[28][197] = 16'h0000;
	mel_filter_coefs[28][198] = 16'h0000;
	mel_filter_coefs[28][199] = 16'h0000;
	mel_filter_coefs[28][200] = 16'h0000;
	mel_filter_coefs[28][201] = 16'h0000;
	mel_filter_coefs[28][202] = 16'h0000;
	mel_filter_coefs[28][203] = 16'h0000;
	mel_filter_coefs[28][204] = 16'h0000;
	mel_filter_coefs[28][205] = 16'h0000;
	mel_filter_coefs[28][206] = 16'h0000;
	mel_filter_coefs[28][207] = 16'h0000;
	mel_filter_coefs[28][208] = 16'h0000;
	mel_filter_coefs[28][209] = 16'h0000;
	mel_filter_coefs[28][210] = 16'h0000;
	mel_filter_coefs[28][211] = 16'h0000;
	mel_filter_coefs[28][212] = 16'h0000;
	mel_filter_coefs[28][213] = 16'h0000;
	mel_filter_coefs[28][214] = 16'h0000;
	mel_filter_coefs[28][215] = 16'h0000;
	mel_filter_coefs[28][216] = 16'h0000;
	mel_filter_coefs[28][217] = 16'h0000;
	mel_filter_coefs[28][218] = 16'h0000;
	mel_filter_coefs[28][219] = 16'h0000;
	mel_filter_coefs[28][220] = 16'h0000;
	mel_filter_coefs[28][221] = 16'h0000;
	mel_filter_coefs[28][222] = 16'h0000;
	mel_filter_coefs[28][223] = 16'h0000;
	mel_filter_coefs[28][224] = 16'h0000;
	mel_filter_coefs[28][225] = 16'h0000;
	mel_filter_coefs[28][226] = 16'h0000;
	mel_filter_coefs[28][227] = 16'h0000;
	mel_filter_coefs[28][228] = 16'h0000;
	mel_filter_coefs[28][229] = 16'h0000;
	mel_filter_coefs[28][230] = 16'h0000;
	mel_filter_coefs[28][231] = 16'h0000;
	mel_filter_coefs[28][232] = 16'h0000;
	mel_filter_coefs[28][233] = 16'h0000;
	mel_filter_coefs[28][234] = 16'h0000;
	mel_filter_coefs[28][235] = 16'h0000;
	mel_filter_coefs[28][236] = 16'h0000;
	mel_filter_coefs[28][237] = 16'h0000;
	mel_filter_coefs[28][238] = 16'h0000;
	mel_filter_coefs[28][239] = 16'h0000;
	mel_filter_coefs[28][240] = 16'h0000;
	mel_filter_coefs[28][241] = 16'h0000;
	mel_filter_coefs[28][242] = 16'h0000;
	mel_filter_coefs[28][243] = 16'h0000;
	mel_filter_coefs[28][244] = 16'h0000;
	mel_filter_coefs[28][245] = 16'h0000;
	mel_filter_coefs[28][246] = 16'h0000;
	mel_filter_coefs[28][247] = 16'h0000;
	mel_filter_coefs[28][248] = 16'h0000;
	mel_filter_coefs[28][249] = 16'h0000;
	mel_filter_coefs[28][250] = 16'h0000;
	mel_filter_coefs[28][251] = 16'h0000;
	mel_filter_coefs[28][252] = 16'h0000;
	mel_filter_coefs[28][253] = 16'h0000;
	mel_filter_coefs[28][254] = 16'h0000;
	mel_filter_coefs[28][255] = 16'h0000;
	mel_filter_coefs[29][0] = 16'h0000;
	mel_filter_coefs[29][1] = 16'h0000;
	mel_filter_coefs[29][2] = 16'h0000;
	mel_filter_coefs[29][3] = 16'h0000;
	mel_filter_coefs[29][4] = 16'h0000;
	mel_filter_coefs[29][5] = 16'h0000;
	mel_filter_coefs[29][6] = 16'h0000;
	mel_filter_coefs[29][7] = 16'h0000;
	mel_filter_coefs[29][8] = 16'h0000;
	mel_filter_coefs[29][9] = 16'h0000;
	mel_filter_coefs[29][10] = 16'h0000;
	mel_filter_coefs[29][11] = 16'h0000;
	mel_filter_coefs[29][12] = 16'h0000;
	mel_filter_coefs[29][13] = 16'h0000;
	mel_filter_coefs[29][14] = 16'h0000;
	mel_filter_coefs[29][15] = 16'h0000;
	mel_filter_coefs[29][16] = 16'h0000;
	mel_filter_coefs[29][17] = 16'h0000;
	mel_filter_coefs[29][18] = 16'h0000;
	mel_filter_coefs[29][19] = 16'h0000;
	mel_filter_coefs[29][20] = 16'h0000;
	mel_filter_coefs[29][21] = 16'h0000;
	mel_filter_coefs[29][22] = 16'h0000;
	mel_filter_coefs[29][23] = 16'h0000;
	mel_filter_coefs[29][24] = 16'h0000;
	mel_filter_coefs[29][25] = 16'h0000;
	mel_filter_coefs[29][26] = 16'h0000;
	mel_filter_coefs[29][27] = 16'h0000;
	mel_filter_coefs[29][28] = 16'h0000;
	mel_filter_coefs[29][29] = 16'h0000;
	mel_filter_coefs[29][30] = 16'h0000;
	mel_filter_coefs[29][31] = 16'h0000;
	mel_filter_coefs[29][32] = 16'h0000;
	mel_filter_coefs[29][33] = 16'h0000;
	mel_filter_coefs[29][34] = 16'h0000;
	mel_filter_coefs[29][35] = 16'h0000;
	mel_filter_coefs[29][36] = 16'h0000;
	mel_filter_coefs[29][37] = 16'h0000;
	mel_filter_coefs[29][38] = 16'h0000;
	mel_filter_coefs[29][39] = 16'h0000;
	mel_filter_coefs[29][40] = 16'h0000;
	mel_filter_coefs[29][41] = 16'h0000;
	mel_filter_coefs[29][42] = 16'h0000;
	mel_filter_coefs[29][43] = 16'h0000;
	mel_filter_coefs[29][44] = 16'h0000;
	mel_filter_coefs[29][45] = 16'h0000;
	mel_filter_coefs[29][46] = 16'h0000;
	mel_filter_coefs[29][47] = 16'h0000;
	mel_filter_coefs[29][48] = 16'h0000;
	mel_filter_coefs[29][49] = 16'h0000;
	mel_filter_coefs[29][50] = 16'h0000;
	mel_filter_coefs[29][51] = 16'h0000;
	mel_filter_coefs[29][52] = 16'h0000;
	mel_filter_coefs[29][53] = 16'h0000;
	mel_filter_coefs[29][54] = 16'h0000;
	mel_filter_coefs[29][55] = 16'h0000;
	mel_filter_coefs[29][56] = 16'h0000;
	mel_filter_coefs[29][57] = 16'h0000;
	mel_filter_coefs[29][58] = 16'h0000;
	mel_filter_coefs[29][59] = 16'h0000;
	mel_filter_coefs[29][60] = 16'h0000;
	mel_filter_coefs[29][61] = 16'h0000;
	mel_filter_coefs[29][62] = 16'h0000;
	mel_filter_coefs[29][63] = 16'h0000;
	mel_filter_coefs[29][64] = 16'h0000;
	mel_filter_coefs[29][65] = 16'h0000;
	mel_filter_coefs[29][66] = 16'h0000;
	mel_filter_coefs[29][67] = 16'h0000;
	mel_filter_coefs[29][68] = 16'h0000;
	mel_filter_coefs[29][69] = 16'h0000;
	mel_filter_coefs[29][70] = 16'h0000;
	mel_filter_coefs[29][71] = 16'h0000;
	mel_filter_coefs[29][72] = 16'h0000;
	mel_filter_coefs[29][73] = 16'h0000;
	mel_filter_coefs[29][74] = 16'h0000;
	mel_filter_coefs[29][75] = 16'h0000;
	mel_filter_coefs[29][76] = 16'h0000;
	mel_filter_coefs[29][77] = 16'h0000;
	mel_filter_coefs[29][78] = 16'h0000;
	mel_filter_coefs[29][79] = 16'h0000;
	mel_filter_coefs[29][80] = 16'h0000;
	mel_filter_coefs[29][81] = 16'h0000;
	mel_filter_coefs[29][82] = 16'h0000;
	mel_filter_coefs[29][83] = 16'h0000;
	mel_filter_coefs[29][84] = 16'h0000;
	mel_filter_coefs[29][85] = 16'h0000;
	mel_filter_coefs[29][86] = 16'h0000;
	mel_filter_coefs[29][87] = 16'h0000;
	mel_filter_coefs[29][88] = 16'h0000;
	mel_filter_coefs[29][89] = 16'h0000;
	mel_filter_coefs[29][90] = 16'h0000;
	mel_filter_coefs[29][91] = 16'h0000;
	mel_filter_coefs[29][92] = 16'h0000;
	mel_filter_coefs[29][93] = 16'h0000;
	mel_filter_coefs[29][94] = 16'h0000;
	mel_filter_coefs[29][95] = 16'h0000;
	mel_filter_coefs[29][96] = 16'h0000;
	mel_filter_coefs[29][97] = 16'h0000;
	mel_filter_coefs[29][98] = 16'h0000;
	mel_filter_coefs[29][99] = 16'h0000;
	mel_filter_coefs[29][100] = 16'h0000;
	mel_filter_coefs[29][101] = 16'h0000;
	mel_filter_coefs[29][102] = 16'h0000;
	mel_filter_coefs[29][103] = 16'h0000;
	mel_filter_coefs[29][104] = 16'h0000;
	mel_filter_coefs[29][105] = 16'h0000;
	mel_filter_coefs[29][106] = 16'h0000;
	mel_filter_coefs[29][107] = 16'h0000;
	mel_filter_coefs[29][108] = 16'h0000;
	mel_filter_coefs[29][109] = 16'h0000;
	mel_filter_coefs[29][110] = 16'h0000;
	mel_filter_coefs[29][111] = 16'h0A59;
	mel_filter_coefs[29][112] = 16'h1992;
	mel_filter_coefs[29][113] = 16'h28CC;
	mel_filter_coefs[29][114] = 16'h3805;
	mel_filter_coefs[29][115] = 16'h473E;
	mel_filter_coefs[29][116] = 16'h5678;
	mel_filter_coefs[29][117] = 16'h65B1;
	mel_filter_coefs[29][118] = 16'h74EA;
	mel_filter_coefs[29][119] = 16'h7C1C;
	mel_filter_coefs[29][120] = 16'h6DCB;
	mel_filter_coefs[29][121] = 16'h5F7A;
	mel_filter_coefs[29][122] = 16'h5129;
	mel_filter_coefs[29][123] = 16'h42D8;
	mel_filter_coefs[29][124] = 16'h3487;
	mel_filter_coefs[29][125] = 16'h2636;
	mel_filter_coefs[29][126] = 16'h17E5;
	mel_filter_coefs[29][127] = 16'h0994;
	mel_filter_coefs[29][128] = 16'h0000;
	mel_filter_coefs[29][129] = 16'h0000;
	mel_filter_coefs[29][130] = 16'h0000;
	mel_filter_coefs[29][131] = 16'h0000;
	mel_filter_coefs[29][132] = 16'h0000;
	mel_filter_coefs[29][133] = 16'h0000;
	mel_filter_coefs[29][134] = 16'h0000;
	mel_filter_coefs[29][135] = 16'h0000;
	mel_filter_coefs[29][136] = 16'h0000;
	mel_filter_coefs[29][137] = 16'h0000;
	mel_filter_coefs[29][138] = 16'h0000;
	mel_filter_coefs[29][139] = 16'h0000;
	mel_filter_coefs[29][140] = 16'h0000;
	mel_filter_coefs[29][141] = 16'h0000;
	mel_filter_coefs[29][142] = 16'h0000;
	mel_filter_coefs[29][143] = 16'h0000;
	mel_filter_coefs[29][144] = 16'h0000;
	mel_filter_coefs[29][145] = 16'h0000;
	mel_filter_coefs[29][146] = 16'h0000;
	mel_filter_coefs[29][147] = 16'h0000;
	mel_filter_coefs[29][148] = 16'h0000;
	mel_filter_coefs[29][149] = 16'h0000;
	mel_filter_coefs[29][150] = 16'h0000;
	mel_filter_coefs[29][151] = 16'h0000;
	mel_filter_coefs[29][152] = 16'h0000;
	mel_filter_coefs[29][153] = 16'h0000;
	mel_filter_coefs[29][154] = 16'h0000;
	mel_filter_coefs[29][155] = 16'h0000;
	mel_filter_coefs[29][156] = 16'h0000;
	mel_filter_coefs[29][157] = 16'h0000;
	mel_filter_coefs[29][158] = 16'h0000;
	mel_filter_coefs[29][159] = 16'h0000;
	mel_filter_coefs[29][160] = 16'h0000;
	mel_filter_coefs[29][161] = 16'h0000;
	mel_filter_coefs[29][162] = 16'h0000;
	mel_filter_coefs[29][163] = 16'h0000;
	mel_filter_coefs[29][164] = 16'h0000;
	mel_filter_coefs[29][165] = 16'h0000;
	mel_filter_coefs[29][166] = 16'h0000;
	mel_filter_coefs[29][167] = 16'h0000;
	mel_filter_coefs[29][168] = 16'h0000;
	mel_filter_coefs[29][169] = 16'h0000;
	mel_filter_coefs[29][170] = 16'h0000;
	mel_filter_coefs[29][171] = 16'h0000;
	mel_filter_coefs[29][172] = 16'h0000;
	mel_filter_coefs[29][173] = 16'h0000;
	mel_filter_coefs[29][174] = 16'h0000;
	mel_filter_coefs[29][175] = 16'h0000;
	mel_filter_coefs[29][176] = 16'h0000;
	mel_filter_coefs[29][177] = 16'h0000;
	mel_filter_coefs[29][178] = 16'h0000;
	mel_filter_coefs[29][179] = 16'h0000;
	mel_filter_coefs[29][180] = 16'h0000;
	mel_filter_coefs[29][181] = 16'h0000;
	mel_filter_coefs[29][182] = 16'h0000;
	mel_filter_coefs[29][183] = 16'h0000;
	mel_filter_coefs[29][184] = 16'h0000;
	mel_filter_coefs[29][185] = 16'h0000;
	mel_filter_coefs[29][186] = 16'h0000;
	mel_filter_coefs[29][187] = 16'h0000;
	mel_filter_coefs[29][188] = 16'h0000;
	mel_filter_coefs[29][189] = 16'h0000;
	mel_filter_coefs[29][190] = 16'h0000;
	mel_filter_coefs[29][191] = 16'h0000;
	mel_filter_coefs[29][192] = 16'h0000;
	mel_filter_coefs[29][193] = 16'h0000;
	mel_filter_coefs[29][194] = 16'h0000;
	mel_filter_coefs[29][195] = 16'h0000;
	mel_filter_coefs[29][196] = 16'h0000;
	mel_filter_coefs[29][197] = 16'h0000;
	mel_filter_coefs[29][198] = 16'h0000;
	mel_filter_coefs[29][199] = 16'h0000;
	mel_filter_coefs[29][200] = 16'h0000;
	mel_filter_coefs[29][201] = 16'h0000;
	mel_filter_coefs[29][202] = 16'h0000;
	mel_filter_coefs[29][203] = 16'h0000;
	mel_filter_coefs[29][204] = 16'h0000;
	mel_filter_coefs[29][205] = 16'h0000;
	mel_filter_coefs[29][206] = 16'h0000;
	mel_filter_coefs[29][207] = 16'h0000;
	mel_filter_coefs[29][208] = 16'h0000;
	mel_filter_coefs[29][209] = 16'h0000;
	mel_filter_coefs[29][210] = 16'h0000;
	mel_filter_coefs[29][211] = 16'h0000;
	mel_filter_coefs[29][212] = 16'h0000;
	mel_filter_coefs[29][213] = 16'h0000;
	mel_filter_coefs[29][214] = 16'h0000;
	mel_filter_coefs[29][215] = 16'h0000;
	mel_filter_coefs[29][216] = 16'h0000;
	mel_filter_coefs[29][217] = 16'h0000;
	mel_filter_coefs[29][218] = 16'h0000;
	mel_filter_coefs[29][219] = 16'h0000;
	mel_filter_coefs[29][220] = 16'h0000;
	mel_filter_coefs[29][221] = 16'h0000;
	mel_filter_coefs[29][222] = 16'h0000;
	mel_filter_coefs[29][223] = 16'h0000;
	mel_filter_coefs[29][224] = 16'h0000;
	mel_filter_coefs[29][225] = 16'h0000;
	mel_filter_coefs[29][226] = 16'h0000;
	mel_filter_coefs[29][227] = 16'h0000;
	mel_filter_coefs[29][228] = 16'h0000;
	mel_filter_coefs[29][229] = 16'h0000;
	mel_filter_coefs[29][230] = 16'h0000;
	mel_filter_coefs[29][231] = 16'h0000;
	mel_filter_coefs[29][232] = 16'h0000;
	mel_filter_coefs[29][233] = 16'h0000;
	mel_filter_coefs[29][234] = 16'h0000;
	mel_filter_coefs[29][235] = 16'h0000;
	mel_filter_coefs[29][236] = 16'h0000;
	mel_filter_coefs[29][237] = 16'h0000;
	mel_filter_coefs[29][238] = 16'h0000;
	mel_filter_coefs[29][239] = 16'h0000;
	mel_filter_coefs[29][240] = 16'h0000;
	mel_filter_coefs[29][241] = 16'h0000;
	mel_filter_coefs[29][242] = 16'h0000;
	mel_filter_coefs[29][243] = 16'h0000;
	mel_filter_coefs[29][244] = 16'h0000;
	mel_filter_coefs[29][245] = 16'h0000;
	mel_filter_coefs[29][246] = 16'h0000;
	mel_filter_coefs[29][247] = 16'h0000;
	mel_filter_coefs[29][248] = 16'h0000;
	mel_filter_coefs[29][249] = 16'h0000;
	mel_filter_coefs[29][250] = 16'h0000;
	mel_filter_coefs[29][251] = 16'h0000;
	mel_filter_coefs[29][252] = 16'h0000;
	mel_filter_coefs[29][253] = 16'h0000;
	mel_filter_coefs[29][254] = 16'h0000;
	mel_filter_coefs[29][255] = 16'h0000;
	mel_filter_coefs[30][0] = 16'h0000;
	mel_filter_coefs[30][1] = 16'h0000;
	mel_filter_coefs[30][2] = 16'h0000;
	mel_filter_coefs[30][3] = 16'h0000;
	mel_filter_coefs[30][4] = 16'h0000;
	mel_filter_coefs[30][5] = 16'h0000;
	mel_filter_coefs[30][6] = 16'h0000;
	mel_filter_coefs[30][7] = 16'h0000;
	mel_filter_coefs[30][8] = 16'h0000;
	mel_filter_coefs[30][9] = 16'h0000;
	mel_filter_coefs[30][10] = 16'h0000;
	mel_filter_coefs[30][11] = 16'h0000;
	mel_filter_coefs[30][12] = 16'h0000;
	mel_filter_coefs[30][13] = 16'h0000;
	mel_filter_coefs[30][14] = 16'h0000;
	mel_filter_coefs[30][15] = 16'h0000;
	mel_filter_coefs[30][16] = 16'h0000;
	mel_filter_coefs[30][17] = 16'h0000;
	mel_filter_coefs[30][18] = 16'h0000;
	mel_filter_coefs[30][19] = 16'h0000;
	mel_filter_coefs[30][20] = 16'h0000;
	mel_filter_coefs[30][21] = 16'h0000;
	mel_filter_coefs[30][22] = 16'h0000;
	mel_filter_coefs[30][23] = 16'h0000;
	mel_filter_coefs[30][24] = 16'h0000;
	mel_filter_coefs[30][25] = 16'h0000;
	mel_filter_coefs[30][26] = 16'h0000;
	mel_filter_coefs[30][27] = 16'h0000;
	mel_filter_coefs[30][28] = 16'h0000;
	mel_filter_coefs[30][29] = 16'h0000;
	mel_filter_coefs[30][30] = 16'h0000;
	mel_filter_coefs[30][31] = 16'h0000;
	mel_filter_coefs[30][32] = 16'h0000;
	mel_filter_coefs[30][33] = 16'h0000;
	mel_filter_coefs[30][34] = 16'h0000;
	mel_filter_coefs[30][35] = 16'h0000;
	mel_filter_coefs[30][36] = 16'h0000;
	mel_filter_coefs[30][37] = 16'h0000;
	mel_filter_coefs[30][38] = 16'h0000;
	mel_filter_coefs[30][39] = 16'h0000;
	mel_filter_coefs[30][40] = 16'h0000;
	mel_filter_coefs[30][41] = 16'h0000;
	mel_filter_coefs[30][42] = 16'h0000;
	mel_filter_coefs[30][43] = 16'h0000;
	mel_filter_coefs[30][44] = 16'h0000;
	mel_filter_coefs[30][45] = 16'h0000;
	mel_filter_coefs[30][46] = 16'h0000;
	mel_filter_coefs[30][47] = 16'h0000;
	mel_filter_coefs[30][48] = 16'h0000;
	mel_filter_coefs[30][49] = 16'h0000;
	mel_filter_coefs[30][50] = 16'h0000;
	mel_filter_coefs[30][51] = 16'h0000;
	mel_filter_coefs[30][52] = 16'h0000;
	mel_filter_coefs[30][53] = 16'h0000;
	mel_filter_coefs[30][54] = 16'h0000;
	mel_filter_coefs[30][55] = 16'h0000;
	mel_filter_coefs[30][56] = 16'h0000;
	mel_filter_coefs[30][57] = 16'h0000;
	mel_filter_coefs[30][58] = 16'h0000;
	mel_filter_coefs[30][59] = 16'h0000;
	mel_filter_coefs[30][60] = 16'h0000;
	mel_filter_coefs[30][61] = 16'h0000;
	mel_filter_coefs[30][62] = 16'h0000;
	mel_filter_coefs[30][63] = 16'h0000;
	mel_filter_coefs[30][64] = 16'h0000;
	mel_filter_coefs[30][65] = 16'h0000;
	mel_filter_coefs[30][66] = 16'h0000;
	mel_filter_coefs[30][67] = 16'h0000;
	mel_filter_coefs[30][68] = 16'h0000;
	mel_filter_coefs[30][69] = 16'h0000;
	mel_filter_coefs[30][70] = 16'h0000;
	mel_filter_coefs[30][71] = 16'h0000;
	mel_filter_coefs[30][72] = 16'h0000;
	mel_filter_coefs[30][73] = 16'h0000;
	mel_filter_coefs[30][74] = 16'h0000;
	mel_filter_coefs[30][75] = 16'h0000;
	mel_filter_coefs[30][76] = 16'h0000;
	mel_filter_coefs[30][77] = 16'h0000;
	mel_filter_coefs[30][78] = 16'h0000;
	mel_filter_coefs[30][79] = 16'h0000;
	mel_filter_coefs[30][80] = 16'h0000;
	mel_filter_coefs[30][81] = 16'h0000;
	mel_filter_coefs[30][82] = 16'h0000;
	mel_filter_coefs[30][83] = 16'h0000;
	mel_filter_coefs[30][84] = 16'h0000;
	mel_filter_coefs[30][85] = 16'h0000;
	mel_filter_coefs[30][86] = 16'h0000;
	mel_filter_coefs[30][87] = 16'h0000;
	mel_filter_coefs[30][88] = 16'h0000;
	mel_filter_coefs[30][89] = 16'h0000;
	mel_filter_coefs[30][90] = 16'h0000;
	mel_filter_coefs[30][91] = 16'h0000;
	mel_filter_coefs[30][92] = 16'h0000;
	mel_filter_coefs[30][93] = 16'h0000;
	mel_filter_coefs[30][94] = 16'h0000;
	mel_filter_coefs[30][95] = 16'h0000;
	mel_filter_coefs[30][96] = 16'h0000;
	mel_filter_coefs[30][97] = 16'h0000;
	mel_filter_coefs[30][98] = 16'h0000;
	mel_filter_coefs[30][99] = 16'h0000;
	mel_filter_coefs[30][100] = 16'h0000;
	mel_filter_coefs[30][101] = 16'h0000;
	mel_filter_coefs[30][102] = 16'h0000;
	mel_filter_coefs[30][103] = 16'h0000;
	mel_filter_coefs[30][104] = 16'h0000;
	mel_filter_coefs[30][105] = 16'h0000;
	mel_filter_coefs[30][106] = 16'h0000;
	mel_filter_coefs[30][107] = 16'h0000;
	mel_filter_coefs[30][108] = 16'h0000;
	mel_filter_coefs[30][109] = 16'h0000;
	mel_filter_coefs[30][110] = 16'h0000;
	mel_filter_coefs[30][111] = 16'h0000;
	mel_filter_coefs[30][112] = 16'h0000;
	mel_filter_coefs[30][113] = 16'h0000;
	mel_filter_coefs[30][114] = 16'h0000;
	mel_filter_coefs[30][115] = 16'h0000;
	mel_filter_coefs[30][116] = 16'h0000;
	mel_filter_coefs[30][117] = 16'h0000;
	mel_filter_coefs[30][118] = 16'h0000;
	mel_filter_coefs[30][119] = 16'h03E4;
	mel_filter_coefs[30][120] = 16'h1235;
	mel_filter_coefs[30][121] = 16'h2086;
	mel_filter_coefs[30][122] = 16'h2ED7;
	mel_filter_coefs[30][123] = 16'h3D28;
	mel_filter_coefs[30][124] = 16'h4B79;
	mel_filter_coefs[30][125] = 16'h59CA;
	mel_filter_coefs[30][126] = 16'h681B;
	mel_filter_coefs[30][127] = 16'h766C;
	mel_filter_coefs[30][128] = 16'h7B8B;
	mel_filter_coefs[30][129] = 16'h6E14;
	mel_filter_coefs[30][130] = 16'h609E;
	mel_filter_coefs[30][131] = 16'h5327;
	mel_filter_coefs[30][132] = 16'h45B1;
	mel_filter_coefs[30][133] = 16'h383A;
	mel_filter_coefs[30][134] = 16'h2AC4;
	mel_filter_coefs[30][135] = 16'h1D4D;
	mel_filter_coefs[30][136] = 16'h0FD7;
	mel_filter_coefs[30][137] = 16'h0260;
	mel_filter_coefs[30][138] = 16'h0000;
	mel_filter_coefs[30][139] = 16'h0000;
	mel_filter_coefs[30][140] = 16'h0000;
	mel_filter_coefs[30][141] = 16'h0000;
	mel_filter_coefs[30][142] = 16'h0000;
	mel_filter_coefs[30][143] = 16'h0000;
	mel_filter_coefs[30][144] = 16'h0000;
	mel_filter_coefs[30][145] = 16'h0000;
	mel_filter_coefs[30][146] = 16'h0000;
	mel_filter_coefs[30][147] = 16'h0000;
	mel_filter_coefs[30][148] = 16'h0000;
	mel_filter_coefs[30][149] = 16'h0000;
	mel_filter_coefs[30][150] = 16'h0000;
	mel_filter_coefs[30][151] = 16'h0000;
	mel_filter_coefs[30][152] = 16'h0000;
	mel_filter_coefs[30][153] = 16'h0000;
	mel_filter_coefs[30][154] = 16'h0000;
	mel_filter_coefs[30][155] = 16'h0000;
	mel_filter_coefs[30][156] = 16'h0000;
	mel_filter_coefs[30][157] = 16'h0000;
	mel_filter_coefs[30][158] = 16'h0000;
	mel_filter_coefs[30][159] = 16'h0000;
	mel_filter_coefs[30][160] = 16'h0000;
	mel_filter_coefs[30][161] = 16'h0000;
	mel_filter_coefs[30][162] = 16'h0000;
	mel_filter_coefs[30][163] = 16'h0000;
	mel_filter_coefs[30][164] = 16'h0000;
	mel_filter_coefs[30][165] = 16'h0000;
	mel_filter_coefs[30][166] = 16'h0000;
	mel_filter_coefs[30][167] = 16'h0000;
	mel_filter_coefs[30][168] = 16'h0000;
	mel_filter_coefs[30][169] = 16'h0000;
	mel_filter_coefs[30][170] = 16'h0000;
	mel_filter_coefs[30][171] = 16'h0000;
	mel_filter_coefs[30][172] = 16'h0000;
	mel_filter_coefs[30][173] = 16'h0000;
	mel_filter_coefs[30][174] = 16'h0000;
	mel_filter_coefs[30][175] = 16'h0000;
	mel_filter_coefs[30][176] = 16'h0000;
	mel_filter_coefs[30][177] = 16'h0000;
	mel_filter_coefs[30][178] = 16'h0000;
	mel_filter_coefs[30][179] = 16'h0000;
	mel_filter_coefs[30][180] = 16'h0000;
	mel_filter_coefs[30][181] = 16'h0000;
	mel_filter_coefs[30][182] = 16'h0000;
	mel_filter_coefs[30][183] = 16'h0000;
	mel_filter_coefs[30][184] = 16'h0000;
	mel_filter_coefs[30][185] = 16'h0000;
	mel_filter_coefs[30][186] = 16'h0000;
	mel_filter_coefs[30][187] = 16'h0000;
	mel_filter_coefs[30][188] = 16'h0000;
	mel_filter_coefs[30][189] = 16'h0000;
	mel_filter_coefs[30][190] = 16'h0000;
	mel_filter_coefs[30][191] = 16'h0000;
	mel_filter_coefs[30][192] = 16'h0000;
	mel_filter_coefs[30][193] = 16'h0000;
	mel_filter_coefs[30][194] = 16'h0000;
	mel_filter_coefs[30][195] = 16'h0000;
	mel_filter_coefs[30][196] = 16'h0000;
	mel_filter_coefs[30][197] = 16'h0000;
	mel_filter_coefs[30][198] = 16'h0000;
	mel_filter_coefs[30][199] = 16'h0000;
	mel_filter_coefs[30][200] = 16'h0000;
	mel_filter_coefs[30][201] = 16'h0000;
	mel_filter_coefs[30][202] = 16'h0000;
	mel_filter_coefs[30][203] = 16'h0000;
	mel_filter_coefs[30][204] = 16'h0000;
	mel_filter_coefs[30][205] = 16'h0000;
	mel_filter_coefs[30][206] = 16'h0000;
	mel_filter_coefs[30][207] = 16'h0000;
	mel_filter_coefs[30][208] = 16'h0000;
	mel_filter_coefs[30][209] = 16'h0000;
	mel_filter_coefs[30][210] = 16'h0000;
	mel_filter_coefs[30][211] = 16'h0000;
	mel_filter_coefs[30][212] = 16'h0000;
	mel_filter_coefs[30][213] = 16'h0000;
	mel_filter_coefs[30][214] = 16'h0000;
	mel_filter_coefs[30][215] = 16'h0000;
	mel_filter_coefs[30][216] = 16'h0000;
	mel_filter_coefs[30][217] = 16'h0000;
	mel_filter_coefs[30][218] = 16'h0000;
	mel_filter_coefs[30][219] = 16'h0000;
	mel_filter_coefs[30][220] = 16'h0000;
	mel_filter_coefs[30][221] = 16'h0000;
	mel_filter_coefs[30][222] = 16'h0000;
	mel_filter_coefs[30][223] = 16'h0000;
	mel_filter_coefs[30][224] = 16'h0000;
	mel_filter_coefs[30][225] = 16'h0000;
	mel_filter_coefs[30][226] = 16'h0000;
	mel_filter_coefs[30][227] = 16'h0000;
	mel_filter_coefs[30][228] = 16'h0000;
	mel_filter_coefs[30][229] = 16'h0000;
	mel_filter_coefs[30][230] = 16'h0000;
	mel_filter_coefs[30][231] = 16'h0000;
	mel_filter_coefs[30][232] = 16'h0000;
	mel_filter_coefs[30][233] = 16'h0000;
	mel_filter_coefs[30][234] = 16'h0000;
	mel_filter_coefs[30][235] = 16'h0000;
	mel_filter_coefs[30][236] = 16'h0000;
	mel_filter_coefs[30][237] = 16'h0000;
	mel_filter_coefs[30][238] = 16'h0000;
	mel_filter_coefs[30][239] = 16'h0000;
	mel_filter_coefs[30][240] = 16'h0000;
	mel_filter_coefs[30][241] = 16'h0000;
	mel_filter_coefs[30][242] = 16'h0000;
	mel_filter_coefs[30][243] = 16'h0000;
	mel_filter_coefs[30][244] = 16'h0000;
	mel_filter_coefs[30][245] = 16'h0000;
	mel_filter_coefs[30][246] = 16'h0000;
	mel_filter_coefs[30][247] = 16'h0000;
	mel_filter_coefs[30][248] = 16'h0000;
	mel_filter_coefs[30][249] = 16'h0000;
	mel_filter_coefs[30][250] = 16'h0000;
	mel_filter_coefs[30][251] = 16'h0000;
	mel_filter_coefs[30][252] = 16'h0000;
	mel_filter_coefs[30][253] = 16'h0000;
	mel_filter_coefs[30][254] = 16'h0000;
	mel_filter_coefs[30][255] = 16'h0000;
	mel_filter_coefs[31][0] = 16'h0000;
	mel_filter_coefs[31][1] = 16'h0000;
	mel_filter_coefs[31][2] = 16'h0000;
	mel_filter_coefs[31][3] = 16'h0000;
	mel_filter_coefs[31][4] = 16'h0000;
	mel_filter_coefs[31][5] = 16'h0000;
	mel_filter_coefs[31][6] = 16'h0000;
	mel_filter_coefs[31][7] = 16'h0000;
	mel_filter_coefs[31][8] = 16'h0000;
	mel_filter_coefs[31][9] = 16'h0000;
	mel_filter_coefs[31][10] = 16'h0000;
	mel_filter_coefs[31][11] = 16'h0000;
	mel_filter_coefs[31][12] = 16'h0000;
	mel_filter_coefs[31][13] = 16'h0000;
	mel_filter_coefs[31][14] = 16'h0000;
	mel_filter_coefs[31][15] = 16'h0000;
	mel_filter_coefs[31][16] = 16'h0000;
	mel_filter_coefs[31][17] = 16'h0000;
	mel_filter_coefs[31][18] = 16'h0000;
	mel_filter_coefs[31][19] = 16'h0000;
	mel_filter_coefs[31][20] = 16'h0000;
	mel_filter_coefs[31][21] = 16'h0000;
	mel_filter_coefs[31][22] = 16'h0000;
	mel_filter_coefs[31][23] = 16'h0000;
	mel_filter_coefs[31][24] = 16'h0000;
	mel_filter_coefs[31][25] = 16'h0000;
	mel_filter_coefs[31][26] = 16'h0000;
	mel_filter_coefs[31][27] = 16'h0000;
	mel_filter_coefs[31][28] = 16'h0000;
	mel_filter_coefs[31][29] = 16'h0000;
	mel_filter_coefs[31][30] = 16'h0000;
	mel_filter_coefs[31][31] = 16'h0000;
	mel_filter_coefs[31][32] = 16'h0000;
	mel_filter_coefs[31][33] = 16'h0000;
	mel_filter_coefs[31][34] = 16'h0000;
	mel_filter_coefs[31][35] = 16'h0000;
	mel_filter_coefs[31][36] = 16'h0000;
	mel_filter_coefs[31][37] = 16'h0000;
	mel_filter_coefs[31][38] = 16'h0000;
	mel_filter_coefs[31][39] = 16'h0000;
	mel_filter_coefs[31][40] = 16'h0000;
	mel_filter_coefs[31][41] = 16'h0000;
	mel_filter_coefs[31][42] = 16'h0000;
	mel_filter_coefs[31][43] = 16'h0000;
	mel_filter_coefs[31][44] = 16'h0000;
	mel_filter_coefs[31][45] = 16'h0000;
	mel_filter_coefs[31][46] = 16'h0000;
	mel_filter_coefs[31][47] = 16'h0000;
	mel_filter_coefs[31][48] = 16'h0000;
	mel_filter_coefs[31][49] = 16'h0000;
	mel_filter_coefs[31][50] = 16'h0000;
	mel_filter_coefs[31][51] = 16'h0000;
	mel_filter_coefs[31][52] = 16'h0000;
	mel_filter_coefs[31][53] = 16'h0000;
	mel_filter_coefs[31][54] = 16'h0000;
	mel_filter_coefs[31][55] = 16'h0000;
	mel_filter_coefs[31][56] = 16'h0000;
	mel_filter_coefs[31][57] = 16'h0000;
	mel_filter_coefs[31][58] = 16'h0000;
	mel_filter_coefs[31][59] = 16'h0000;
	mel_filter_coefs[31][60] = 16'h0000;
	mel_filter_coefs[31][61] = 16'h0000;
	mel_filter_coefs[31][62] = 16'h0000;
	mel_filter_coefs[31][63] = 16'h0000;
	mel_filter_coefs[31][64] = 16'h0000;
	mel_filter_coefs[31][65] = 16'h0000;
	mel_filter_coefs[31][66] = 16'h0000;
	mel_filter_coefs[31][67] = 16'h0000;
	mel_filter_coefs[31][68] = 16'h0000;
	mel_filter_coefs[31][69] = 16'h0000;
	mel_filter_coefs[31][70] = 16'h0000;
	mel_filter_coefs[31][71] = 16'h0000;
	mel_filter_coefs[31][72] = 16'h0000;
	mel_filter_coefs[31][73] = 16'h0000;
	mel_filter_coefs[31][74] = 16'h0000;
	mel_filter_coefs[31][75] = 16'h0000;
	mel_filter_coefs[31][76] = 16'h0000;
	mel_filter_coefs[31][77] = 16'h0000;
	mel_filter_coefs[31][78] = 16'h0000;
	mel_filter_coefs[31][79] = 16'h0000;
	mel_filter_coefs[31][80] = 16'h0000;
	mel_filter_coefs[31][81] = 16'h0000;
	mel_filter_coefs[31][82] = 16'h0000;
	mel_filter_coefs[31][83] = 16'h0000;
	mel_filter_coefs[31][84] = 16'h0000;
	mel_filter_coefs[31][85] = 16'h0000;
	mel_filter_coefs[31][86] = 16'h0000;
	mel_filter_coefs[31][87] = 16'h0000;
	mel_filter_coefs[31][88] = 16'h0000;
	mel_filter_coefs[31][89] = 16'h0000;
	mel_filter_coefs[31][90] = 16'h0000;
	mel_filter_coefs[31][91] = 16'h0000;
	mel_filter_coefs[31][92] = 16'h0000;
	mel_filter_coefs[31][93] = 16'h0000;
	mel_filter_coefs[31][94] = 16'h0000;
	mel_filter_coefs[31][95] = 16'h0000;
	mel_filter_coefs[31][96] = 16'h0000;
	mel_filter_coefs[31][97] = 16'h0000;
	mel_filter_coefs[31][98] = 16'h0000;
	mel_filter_coefs[31][99] = 16'h0000;
	mel_filter_coefs[31][100] = 16'h0000;
	mel_filter_coefs[31][101] = 16'h0000;
	mel_filter_coefs[31][102] = 16'h0000;
	mel_filter_coefs[31][103] = 16'h0000;
	mel_filter_coefs[31][104] = 16'h0000;
	mel_filter_coefs[31][105] = 16'h0000;
	mel_filter_coefs[31][106] = 16'h0000;
	mel_filter_coefs[31][107] = 16'h0000;
	mel_filter_coefs[31][108] = 16'h0000;
	mel_filter_coefs[31][109] = 16'h0000;
	mel_filter_coefs[31][110] = 16'h0000;
	mel_filter_coefs[31][111] = 16'h0000;
	mel_filter_coefs[31][112] = 16'h0000;
	mel_filter_coefs[31][113] = 16'h0000;
	mel_filter_coefs[31][114] = 16'h0000;
	mel_filter_coefs[31][115] = 16'h0000;
	mel_filter_coefs[31][116] = 16'h0000;
	mel_filter_coefs[31][117] = 16'h0000;
	mel_filter_coefs[31][118] = 16'h0000;
	mel_filter_coefs[31][119] = 16'h0000;
	mel_filter_coefs[31][120] = 16'h0000;
	mel_filter_coefs[31][121] = 16'h0000;
	mel_filter_coefs[31][122] = 16'h0000;
	mel_filter_coefs[31][123] = 16'h0000;
	mel_filter_coefs[31][124] = 16'h0000;
	mel_filter_coefs[31][125] = 16'h0000;
	mel_filter_coefs[31][126] = 16'h0000;
	mel_filter_coefs[31][127] = 16'h0000;
	mel_filter_coefs[31][128] = 16'h0475;
	mel_filter_coefs[31][129] = 16'h11EC;
	mel_filter_coefs[31][130] = 16'h1F62;
	mel_filter_coefs[31][131] = 16'h2CD9;
	mel_filter_coefs[31][132] = 16'h3A4F;
	mel_filter_coefs[31][133] = 16'h47C6;
	mel_filter_coefs[31][134] = 16'h553C;
	mel_filter_coefs[31][135] = 16'h62B3;
	mel_filter_coefs[31][136] = 16'h7029;
	mel_filter_coefs[31][137] = 16'h7DA0;
	mel_filter_coefs[31][138] = 16'h7593;
	mel_filter_coefs[31][139] = 16'h68EA;
	mel_filter_coefs[31][140] = 16'h5C41;
	mel_filter_coefs[31][141] = 16'h4F98;
	mel_filter_coefs[31][142] = 16'h42EF;
	mel_filter_coefs[31][143] = 16'h3646;
	mel_filter_coefs[31][144] = 16'h299C;
	mel_filter_coefs[31][145] = 16'h1CF3;
	mel_filter_coefs[31][146] = 16'h104A;
	mel_filter_coefs[31][147] = 16'h03A1;
	mel_filter_coefs[31][148] = 16'h0000;
	mel_filter_coefs[31][149] = 16'h0000;
	mel_filter_coefs[31][150] = 16'h0000;
	mel_filter_coefs[31][151] = 16'h0000;
	mel_filter_coefs[31][152] = 16'h0000;
	mel_filter_coefs[31][153] = 16'h0000;
	mel_filter_coefs[31][154] = 16'h0000;
	mel_filter_coefs[31][155] = 16'h0000;
	mel_filter_coefs[31][156] = 16'h0000;
	mel_filter_coefs[31][157] = 16'h0000;
	mel_filter_coefs[31][158] = 16'h0000;
	mel_filter_coefs[31][159] = 16'h0000;
	mel_filter_coefs[31][160] = 16'h0000;
	mel_filter_coefs[31][161] = 16'h0000;
	mel_filter_coefs[31][162] = 16'h0000;
	mel_filter_coefs[31][163] = 16'h0000;
	mel_filter_coefs[31][164] = 16'h0000;
	mel_filter_coefs[31][165] = 16'h0000;
	mel_filter_coefs[31][166] = 16'h0000;
	mel_filter_coefs[31][167] = 16'h0000;
	mel_filter_coefs[31][168] = 16'h0000;
	mel_filter_coefs[31][169] = 16'h0000;
	mel_filter_coefs[31][170] = 16'h0000;
	mel_filter_coefs[31][171] = 16'h0000;
	mel_filter_coefs[31][172] = 16'h0000;
	mel_filter_coefs[31][173] = 16'h0000;
	mel_filter_coefs[31][174] = 16'h0000;
	mel_filter_coefs[31][175] = 16'h0000;
	mel_filter_coefs[31][176] = 16'h0000;
	mel_filter_coefs[31][177] = 16'h0000;
	mel_filter_coefs[31][178] = 16'h0000;
	mel_filter_coefs[31][179] = 16'h0000;
	mel_filter_coefs[31][180] = 16'h0000;
	mel_filter_coefs[31][181] = 16'h0000;
	mel_filter_coefs[31][182] = 16'h0000;
	mel_filter_coefs[31][183] = 16'h0000;
	mel_filter_coefs[31][184] = 16'h0000;
	mel_filter_coefs[31][185] = 16'h0000;
	mel_filter_coefs[31][186] = 16'h0000;
	mel_filter_coefs[31][187] = 16'h0000;
	mel_filter_coefs[31][188] = 16'h0000;
	mel_filter_coefs[31][189] = 16'h0000;
	mel_filter_coefs[31][190] = 16'h0000;
	mel_filter_coefs[31][191] = 16'h0000;
	mel_filter_coefs[31][192] = 16'h0000;
	mel_filter_coefs[31][193] = 16'h0000;
	mel_filter_coefs[31][194] = 16'h0000;
	mel_filter_coefs[31][195] = 16'h0000;
	mel_filter_coefs[31][196] = 16'h0000;
	mel_filter_coefs[31][197] = 16'h0000;
	mel_filter_coefs[31][198] = 16'h0000;
	mel_filter_coefs[31][199] = 16'h0000;
	mel_filter_coefs[31][200] = 16'h0000;
	mel_filter_coefs[31][201] = 16'h0000;
	mel_filter_coefs[31][202] = 16'h0000;
	mel_filter_coefs[31][203] = 16'h0000;
	mel_filter_coefs[31][204] = 16'h0000;
	mel_filter_coefs[31][205] = 16'h0000;
	mel_filter_coefs[31][206] = 16'h0000;
	mel_filter_coefs[31][207] = 16'h0000;
	mel_filter_coefs[31][208] = 16'h0000;
	mel_filter_coefs[31][209] = 16'h0000;
	mel_filter_coefs[31][210] = 16'h0000;
	mel_filter_coefs[31][211] = 16'h0000;
	mel_filter_coefs[31][212] = 16'h0000;
	mel_filter_coefs[31][213] = 16'h0000;
	mel_filter_coefs[31][214] = 16'h0000;
	mel_filter_coefs[31][215] = 16'h0000;
	mel_filter_coefs[31][216] = 16'h0000;
	mel_filter_coefs[31][217] = 16'h0000;
	mel_filter_coefs[31][218] = 16'h0000;
	mel_filter_coefs[31][219] = 16'h0000;
	mel_filter_coefs[31][220] = 16'h0000;
	mel_filter_coefs[31][221] = 16'h0000;
	mel_filter_coefs[31][222] = 16'h0000;
	mel_filter_coefs[31][223] = 16'h0000;
	mel_filter_coefs[31][224] = 16'h0000;
	mel_filter_coefs[31][225] = 16'h0000;
	mel_filter_coefs[31][226] = 16'h0000;
	mel_filter_coefs[31][227] = 16'h0000;
	mel_filter_coefs[31][228] = 16'h0000;
	mel_filter_coefs[31][229] = 16'h0000;
	mel_filter_coefs[31][230] = 16'h0000;
	mel_filter_coefs[31][231] = 16'h0000;
	mel_filter_coefs[31][232] = 16'h0000;
	mel_filter_coefs[31][233] = 16'h0000;
	mel_filter_coefs[31][234] = 16'h0000;
	mel_filter_coefs[31][235] = 16'h0000;
	mel_filter_coefs[31][236] = 16'h0000;
	mel_filter_coefs[31][237] = 16'h0000;
	mel_filter_coefs[31][238] = 16'h0000;
	mel_filter_coefs[31][239] = 16'h0000;
	mel_filter_coefs[31][240] = 16'h0000;
	mel_filter_coefs[31][241] = 16'h0000;
	mel_filter_coefs[31][242] = 16'h0000;
	mel_filter_coefs[31][243] = 16'h0000;
	mel_filter_coefs[31][244] = 16'h0000;
	mel_filter_coefs[31][245] = 16'h0000;
	mel_filter_coefs[31][246] = 16'h0000;
	mel_filter_coefs[31][247] = 16'h0000;
	mel_filter_coefs[31][248] = 16'h0000;
	mel_filter_coefs[31][249] = 16'h0000;
	mel_filter_coefs[31][250] = 16'h0000;
	mel_filter_coefs[31][251] = 16'h0000;
	mel_filter_coefs[31][252] = 16'h0000;
	mel_filter_coefs[31][253] = 16'h0000;
	mel_filter_coefs[31][254] = 16'h0000;
	mel_filter_coefs[31][255] = 16'h0000;
	mel_filter_coefs[32][0] = 16'h0000;
	mel_filter_coefs[32][1] = 16'h0000;
	mel_filter_coefs[32][2] = 16'h0000;
	mel_filter_coefs[32][3] = 16'h0000;
	mel_filter_coefs[32][4] = 16'h0000;
	mel_filter_coefs[32][5] = 16'h0000;
	mel_filter_coefs[32][6] = 16'h0000;
	mel_filter_coefs[32][7] = 16'h0000;
	mel_filter_coefs[32][8] = 16'h0000;
	mel_filter_coefs[32][9] = 16'h0000;
	mel_filter_coefs[32][10] = 16'h0000;
	mel_filter_coefs[32][11] = 16'h0000;
	mel_filter_coefs[32][12] = 16'h0000;
	mel_filter_coefs[32][13] = 16'h0000;
	mel_filter_coefs[32][14] = 16'h0000;
	mel_filter_coefs[32][15] = 16'h0000;
	mel_filter_coefs[32][16] = 16'h0000;
	mel_filter_coefs[32][17] = 16'h0000;
	mel_filter_coefs[32][18] = 16'h0000;
	mel_filter_coefs[32][19] = 16'h0000;
	mel_filter_coefs[32][20] = 16'h0000;
	mel_filter_coefs[32][21] = 16'h0000;
	mel_filter_coefs[32][22] = 16'h0000;
	mel_filter_coefs[32][23] = 16'h0000;
	mel_filter_coefs[32][24] = 16'h0000;
	mel_filter_coefs[32][25] = 16'h0000;
	mel_filter_coefs[32][26] = 16'h0000;
	mel_filter_coefs[32][27] = 16'h0000;
	mel_filter_coefs[32][28] = 16'h0000;
	mel_filter_coefs[32][29] = 16'h0000;
	mel_filter_coefs[32][30] = 16'h0000;
	mel_filter_coefs[32][31] = 16'h0000;
	mel_filter_coefs[32][32] = 16'h0000;
	mel_filter_coefs[32][33] = 16'h0000;
	mel_filter_coefs[32][34] = 16'h0000;
	mel_filter_coefs[32][35] = 16'h0000;
	mel_filter_coefs[32][36] = 16'h0000;
	mel_filter_coefs[32][37] = 16'h0000;
	mel_filter_coefs[32][38] = 16'h0000;
	mel_filter_coefs[32][39] = 16'h0000;
	mel_filter_coefs[32][40] = 16'h0000;
	mel_filter_coefs[32][41] = 16'h0000;
	mel_filter_coefs[32][42] = 16'h0000;
	mel_filter_coefs[32][43] = 16'h0000;
	mel_filter_coefs[32][44] = 16'h0000;
	mel_filter_coefs[32][45] = 16'h0000;
	mel_filter_coefs[32][46] = 16'h0000;
	mel_filter_coefs[32][47] = 16'h0000;
	mel_filter_coefs[32][48] = 16'h0000;
	mel_filter_coefs[32][49] = 16'h0000;
	mel_filter_coefs[32][50] = 16'h0000;
	mel_filter_coefs[32][51] = 16'h0000;
	mel_filter_coefs[32][52] = 16'h0000;
	mel_filter_coefs[32][53] = 16'h0000;
	mel_filter_coefs[32][54] = 16'h0000;
	mel_filter_coefs[32][55] = 16'h0000;
	mel_filter_coefs[32][56] = 16'h0000;
	mel_filter_coefs[32][57] = 16'h0000;
	mel_filter_coefs[32][58] = 16'h0000;
	mel_filter_coefs[32][59] = 16'h0000;
	mel_filter_coefs[32][60] = 16'h0000;
	mel_filter_coefs[32][61] = 16'h0000;
	mel_filter_coefs[32][62] = 16'h0000;
	mel_filter_coefs[32][63] = 16'h0000;
	mel_filter_coefs[32][64] = 16'h0000;
	mel_filter_coefs[32][65] = 16'h0000;
	mel_filter_coefs[32][66] = 16'h0000;
	mel_filter_coefs[32][67] = 16'h0000;
	mel_filter_coefs[32][68] = 16'h0000;
	mel_filter_coefs[32][69] = 16'h0000;
	mel_filter_coefs[32][70] = 16'h0000;
	mel_filter_coefs[32][71] = 16'h0000;
	mel_filter_coefs[32][72] = 16'h0000;
	mel_filter_coefs[32][73] = 16'h0000;
	mel_filter_coefs[32][74] = 16'h0000;
	mel_filter_coefs[32][75] = 16'h0000;
	mel_filter_coefs[32][76] = 16'h0000;
	mel_filter_coefs[32][77] = 16'h0000;
	mel_filter_coefs[32][78] = 16'h0000;
	mel_filter_coefs[32][79] = 16'h0000;
	mel_filter_coefs[32][80] = 16'h0000;
	mel_filter_coefs[32][81] = 16'h0000;
	mel_filter_coefs[32][82] = 16'h0000;
	mel_filter_coefs[32][83] = 16'h0000;
	mel_filter_coefs[32][84] = 16'h0000;
	mel_filter_coefs[32][85] = 16'h0000;
	mel_filter_coefs[32][86] = 16'h0000;
	mel_filter_coefs[32][87] = 16'h0000;
	mel_filter_coefs[32][88] = 16'h0000;
	mel_filter_coefs[32][89] = 16'h0000;
	mel_filter_coefs[32][90] = 16'h0000;
	mel_filter_coefs[32][91] = 16'h0000;
	mel_filter_coefs[32][92] = 16'h0000;
	mel_filter_coefs[32][93] = 16'h0000;
	mel_filter_coefs[32][94] = 16'h0000;
	mel_filter_coefs[32][95] = 16'h0000;
	mel_filter_coefs[32][96] = 16'h0000;
	mel_filter_coefs[32][97] = 16'h0000;
	mel_filter_coefs[32][98] = 16'h0000;
	mel_filter_coefs[32][99] = 16'h0000;
	mel_filter_coefs[32][100] = 16'h0000;
	mel_filter_coefs[32][101] = 16'h0000;
	mel_filter_coefs[32][102] = 16'h0000;
	mel_filter_coefs[32][103] = 16'h0000;
	mel_filter_coefs[32][104] = 16'h0000;
	mel_filter_coefs[32][105] = 16'h0000;
	mel_filter_coefs[32][106] = 16'h0000;
	mel_filter_coefs[32][107] = 16'h0000;
	mel_filter_coefs[32][108] = 16'h0000;
	mel_filter_coefs[32][109] = 16'h0000;
	mel_filter_coefs[32][110] = 16'h0000;
	mel_filter_coefs[32][111] = 16'h0000;
	mel_filter_coefs[32][112] = 16'h0000;
	mel_filter_coefs[32][113] = 16'h0000;
	mel_filter_coefs[32][114] = 16'h0000;
	mel_filter_coefs[32][115] = 16'h0000;
	mel_filter_coefs[32][116] = 16'h0000;
	mel_filter_coefs[32][117] = 16'h0000;
	mel_filter_coefs[32][118] = 16'h0000;
	mel_filter_coefs[32][119] = 16'h0000;
	mel_filter_coefs[32][120] = 16'h0000;
	mel_filter_coefs[32][121] = 16'h0000;
	mel_filter_coefs[32][122] = 16'h0000;
	mel_filter_coefs[32][123] = 16'h0000;
	mel_filter_coefs[32][124] = 16'h0000;
	mel_filter_coefs[32][125] = 16'h0000;
	mel_filter_coefs[32][126] = 16'h0000;
	mel_filter_coefs[32][127] = 16'h0000;
	mel_filter_coefs[32][128] = 16'h0000;
	mel_filter_coefs[32][129] = 16'h0000;
	mel_filter_coefs[32][130] = 16'h0000;
	mel_filter_coefs[32][131] = 16'h0000;
	mel_filter_coefs[32][132] = 16'h0000;
	mel_filter_coefs[32][133] = 16'h0000;
	mel_filter_coefs[32][134] = 16'h0000;
	mel_filter_coefs[32][135] = 16'h0000;
	mel_filter_coefs[32][136] = 16'h0000;
	mel_filter_coefs[32][137] = 16'h0000;
	mel_filter_coefs[32][138] = 16'h0A6D;
	mel_filter_coefs[32][139] = 16'h1716;
	mel_filter_coefs[32][140] = 16'h23BF;
	mel_filter_coefs[32][141] = 16'h3068;
	mel_filter_coefs[32][142] = 16'h3D11;
	mel_filter_coefs[32][143] = 16'h49BA;
	mel_filter_coefs[32][144] = 16'h5664;
	mel_filter_coefs[32][145] = 16'h630D;
	mel_filter_coefs[32][146] = 16'h6FB6;
	mel_filter_coefs[32][147] = 16'h7C5F;
	mel_filter_coefs[32][148] = 16'h7782;
	mel_filter_coefs[32][149] = 16'h6B9A;
	mel_filter_coefs[32][150] = 16'h5FB2;
	mel_filter_coefs[32][151] = 16'h53CA;
	mel_filter_coefs[32][152] = 16'h47E3;
	mel_filter_coefs[32][153] = 16'h3BFB;
	mel_filter_coefs[32][154] = 16'h3013;
	mel_filter_coefs[32][155] = 16'h242B;
	mel_filter_coefs[32][156] = 16'h1843;
	mel_filter_coefs[32][157] = 16'h0C5B;
	mel_filter_coefs[32][158] = 16'h0073;
	mel_filter_coefs[32][159] = 16'h0000;
	mel_filter_coefs[32][160] = 16'h0000;
	mel_filter_coefs[32][161] = 16'h0000;
	mel_filter_coefs[32][162] = 16'h0000;
	mel_filter_coefs[32][163] = 16'h0000;
	mel_filter_coefs[32][164] = 16'h0000;
	mel_filter_coefs[32][165] = 16'h0000;
	mel_filter_coefs[32][166] = 16'h0000;
	mel_filter_coefs[32][167] = 16'h0000;
	mel_filter_coefs[32][168] = 16'h0000;
	mel_filter_coefs[32][169] = 16'h0000;
	mel_filter_coefs[32][170] = 16'h0000;
	mel_filter_coefs[32][171] = 16'h0000;
	mel_filter_coefs[32][172] = 16'h0000;
	mel_filter_coefs[32][173] = 16'h0000;
	mel_filter_coefs[32][174] = 16'h0000;
	mel_filter_coefs[32][175] = 16'h0000;
	mel_filter_coefs[32][176] = 16'h0000;
	mel_filter_coefs[32][177] = 16'h0000;
	mel_filter_coefs[32][178] = 16'h0000;
	mel_filter_coefs[32][179] = 16'h0000;
	mel_filter_coefs[32][180] = 16'h0000;
	mel_filter_coefs[32][181] = 16'h0000;
	mel_filter_coefs[32][182] = 16'h0000;
	mel_filter_coefs[32][183] = 16'h0000;
	mel_filter_coefs[32][184] = 16'h0000;
	mel_filter_coefs[32][185] = 16'h0000;
	mel_filter_coefs[32][186] = 16'h0000;
	mel_filter_coefs[32][187] = 16'h0000;
	mel_filter_coefs[32][188] = 16'h0000;
	mel_filter_coefs[32][189] = 16'h0000;
	mel_filter_coefs[32][190] = 16'h0000;
	mel_filter_coefs[32][191] = 16'h0000;
	mel_filter_coefs[32][192] = 16'h0000;
	mel_filter_coefs[32][193] = 16'h0000;
	mel_filter_coefs[32][194] = 16'h0000;
	mel_filter_coefs[32][195] = 16'h0000;
	mel_filter_coefs[32][196] = 16'h0000;
	mel_filter_coefs[32][197] = 16'h0000;
	mel_filter_coefs[32][198] = 16'h0000;
	mel_filter_coefs[32][199] = 16'h0000;
	mel_filter_coefs[32][200] = 16'h0000;
	mel_filter_coefs[32][201] = 16'h0000;
	mel_filter_coefs[32][202] = 16'h0000;
	mel_filter_coefs[32][203] = 16'h0000;
	mel_filter_coefs[32][204] = 16'h0000;
	mel_filter_coefs[32][205] = 16'h0000;
	mel_filter_coefs[32][206] = 16'h0000;
	mel_filter_coefs[32][207] = 16'h0000;
	mel_filter_coefs[32][208] = 16'h0000;
	mel_filter_coefs[32][209] = 16'h0000;
	mel_filter_coefs[32][210] = 16'h0000;
	mel_filter_coefs[32][211] = 16'h0000;
	mel_filter_coefs[32][212] = 16'h0000;
	mel_filter_coefs[32][213] = 16'h0000;
	mel_filter_coefs[32][214] = 16'h0000;
	mel_filter_coefs[32][215] = 16'h0000;
	mel_filter_coefs[32][216] = 16'h0000;
	mel_filter_coefs[32][217] = 16'h0000;
	mel_filter_coefs[32][218] = 16'h0000;
	mel_filter_coefs[32][219] = 16'h0000;
	mel_filter_coefs[32][220] = 16'h0000;
	mel_filter_coefs[32][221] = 16'h0000;
	mel_filter_coefs[32][222] = 16'h0000;
	mel_filter_coefs[32][223] = 16'h0000;
	mel_filter_coefs[32][224] = 16'h0000;
	mel_filter_coefs[32][225] = 16'h0000;
	mel_filter_coefs[32][226] = 16'h0000;
	mel_filter_coefs[32][227] = 16'h0000;
	mel_filter_coefs[32][228] = 16'h0000;
	mel_filter_coefs[32][229] = 16'h0000;
	mel_filter_coefs[32][230] = 16'h0000;
	mel_filter_coefs[32][231] = 16'h0000;
	mel_filter_coefs[32][232] = 16'h0000;
	mel_filter_coefs[32][233] = 16'h0000;
	mel_filter_coefs[32][234] = 16'h0000;
	mel_filter_coefs[32][235] = 16'h0000;
	mel_filter_coefs[32][236] = 16'h0000;
	mel_filter_coefs[32][237] = 16'h0000;
	mel_filter_coefs[32][238] = 16'h0000;
	mel_filter_coefs[32][239] = 16'h0000;
	mel_filter_coefs[32][240] = 16'h0000;
	mel_filter_coefs[32][241] = 16'h0000;
	mel_filter_coefs[32][242] = 16'h0000;
	mel_filter_coefs[32][243] = 16'h0000;
	mel_filter_coefs[32][244] = 16'h0000;
	mel_filter_coefs[32][245] = 16'h0000;
	mel_filter_coefs[32][246] = 16'h0000;
	mel_filter_coefs[32][247] = 16'h0000;
	mel_filter_coefs[32][248] = 16'h0000;
	mel_filter_coefs[32][249] = 16'h0000;
	mel_filter_coefs[32][250] = 16'h0000;
	mel_filter_coefs[32][251] = 16'h0000;
	mel_filter_coefs[32][252] = 16'h0000;
	mel_filter_coefs[32][253] = 16'h0000;
	mel_filter_coefs[32][254] = 16'h0000;
	mel_filter_coefs[32][255] = 16'h0000;
	mel_filter_coefs[33][0] = 16'h0000;
	mel_filter_coefs[33][1] = 16'h0000;
	mel_filter_coefs[33][2] = 16'h0000;
	mel_filter_coefs[33][3] = 16'h0000;
	mel_filter_coefs[33][4] = 16'h0000;
	mel_filter_coefs[33][5] = 16'h0000;
	mel_filter_coefs[33][6] = 16'h0000;
	mel_filter_coefs[33][7] = 16'h0000;
	mel_filter_coefs[33][8] = 16'h0000;
	mel_filter_coefs[33][9] = 16'h0000;
	mel_filter_coefs[33][10] = 16'h0000;
	mel_filter_coefs[33][11] = 16'h0000;
	mel_filter_coefs[33][12] = 16'h0000;
	mel_filter_coefs[33][13] = 16'h0000;
	mel_filter_coefs[33][14] = 16'h0000;
	mel_filter_coefs[33][15] = 16'h0000;
	mel_filter_coefs[33][16] = 16'h0000;
	mel_filter_coefs[33][17] = 16'h0000;
	mel_filter_coefs[33][18] = 16'h0000;
	mel_filter_coefs[33][19] = 16'h0000;
	mel_filter_coefs[33][20] = 16'h0000;
	mel_filter_coefs[33][21] = 16'h0000;
	mel_filter_coefs[33][22] = 16'h0000;
	mel_filter_coefs[33][23] = 16'h0000;
	mel_filter_coefs[33][24] = 16'h0000;
	mel_filter_coefs[33][25] = 16'h0000;
	mel_filter_coefs[33][26] = 16'h0000;
	mel_filter_coefs[33][27] = 16'h0000;
	mel_filter_coefs[33][28] = 16'h0000;
	mel_filter_coefs[33][29] = 16'h0000;
	mel_filter_coefs[33][30] = 16'h0000;
	mel_filter_coefs[33][31] = 16'h0000;
	mel_filter_coefs[33][32] = 16'h0000;
	mel_filter_coefs[33][33] = 16'h0000;
	mel_filter_coefs[33][34] = 16'h0000;
	mel_filter_coefs[33][35] = 16'h0000;
	mel_filter_coefs[33][36] = 16'h0000;
	mel_filter_coefs[33][37] = 16'h0000;
	mel_filter_coefs[33][38] = 16'h0000;
	mel_filter_coefs[33][39] = 16'h0000;
	mel_filter_coefs[33][40] = 16'h0000;
	mel_filter_coefs[33][41] = 16'h0000;
	mel_filter_coefs[33][42] = 16'h0000;
	mel_filter_coefs[33][43] = 16'h0000;
	mel_filter_coefs[33][44] = 16'h0000;
	mel_filter_coefs[33][45] = 16'h0000;
	mel_filter_coefs[33][46] = 16'h0000;
	mel_filter_coefs[33][47] = 16'h0000;
	mel_filter_coefs[33][48] = 16'h0000;
	mel_filter_coefs[33][49] = 16'h0000;
	mel_filter_coefs[33][50] = 16'h0000;
	mel_filter_coefs[33][51] = 16'h0000;
	mel_filter_coefs[33][52] = 16'h0000;
	mel_filter_coefs[33][53] = 16'h0000;
	mel_filter_coefs[33][54] = 16'h0000;
	mel_filter_coefs[33][55] = 16'h0000;
	mel_filter_coefs[33][56] = 16'h0000;
	mel_filter_coefs[33][57] = 16'h0000;
	mel_filter_coefs[33][58] = 16'h0000;
	mel_filter_coefs[33][59] = 16'h0000;
	mel_filter_coefs[33][60] = 16'h0000;
	mel_filter_coefs[33][61] = 16'h0000;
	mel_filter_coefs[33][62] = 16'h0000;
	mel_filter_coefs[33][63] = 16'h0000;
	mel_filter_coefs[33][64] = 16'h0000;
	mel_filter_coefs[33][65] = 16'h0000;
	mel_filter_coefs[33][66] = 16'h0000;
	mel_filter_coefs[33][67] = 16'h0000;
	mel_filter_coefs[33][68] = 16'h0000;
	mel_filter_coefs[33][69] = 16'h0000;
	mel_filter_coefs[33][70] = 16'h0000;
	mel_filter_coefs[33][71] = 16'h0000;
	mel_filter_coefs[33][72] = 16'h0000;
	mel_filter_coefs[33][73] = 16'h0000;
	mel_filter_coefs[33][74] = 16'h0000;
	mel_filter_coefs[33][75] = 16'h0000;
	mel_filter_coefs[33][76] = 16'h0000;
	mel_filter_coefs[33][77] = 16'h0000;
	mel_filter_coefs[33][78] = 16'h0000;
	mel_filter_coefs[33][79] = 16'h0000;
	mel_filter_coefs[33][80] = 16'h0000;
	mel_filter_coefs[33][81] = 16'h0000;
	mel_filter_coefs[33][82] = 16'h0000;
	mel_filter_coefs[33][83] = 16'h0000;
	mel_filter_coefs[33][84] = 16'h0000;
	mel_filter_coefs[33][85] = 16'h0000;
	mel_filter_coefs[33][86] = 16'h0000;
	mel_filter_coefs[33][87] = 16'h0000;
	mel_filter_coefs[33][88] = 16'h0000;
	mel_filter_coefs[33][89] = 16'h0000;
	mel_filter_coefs[33][90] = 16'h0000;
	mel_filter_coefs[33][91] = 16'h0000;
	mel_filter_coefs[33][92] = 16'h0000;
	mel_filter_coefs[33][93] = 16'h0000;
	mel_filter_coefs[33][94] = 16'h0000;
	mel_filter_coefs[33][95] = 16'h0000;
	mel_filter_coefs[33][96] = 16'h0000;
	mel_filter_coefs[33][97] = 16'h0000;
	mel_filter_coefs[33][98] = 16'h0000;
	mel_filter_coefs[33][99] = 16'h0000;
	mel_filter_coefs[33][100] = 16'h0000;
	mel_filter_coefs[33][101] = 16'h0000;
	mel_filter_coefs[33][102] = 16'h0000;
	mel_filter_coefs[33][103] = 16'h0000;
	mel_filter_coefs[33][104] = 16'h0000;
	mel_filter_coefs[33][105] = 16'h0000;
	mel_filter_coefs[33][106] = 16'h0000;
	mel_filter_coefs[33][107] = 16'h0000;
	mel_filter_coefs[33][108] = 16'h0000;
	mel_filter_coefs[33][109] = 16'h0000;
	mel_filter_coefs[33][110] = 16'h0000;
	mel_filter_coefs[33][111] = 16'h0000;
	mel_filter_coefs[33][112] = 16'h0000;
	mel_filter_coefs[33][113] = 16'h0000;
	mel_filter_coefs[33][114] = 16'h0000;
	mel_filter_coefs[33][115] = 16'h0000;
	mel_filter_coefs[33][116] = 16'h0000;
	mel_filter_coefs[33][117] = 16'h0000;
	mel_filter_coefs[33][118] = 16'h0000;
	mel_filter_coefs[33][119] = 16'h0000;
	mel_filter_coefs[33][120] = 16'h0000;
	mel_filter_coefs[33][121] = 16'h0000;
	mel_filter_coefs[33][122] = 16'h0000;
	mel_filter_coefs[33][123] = 16'h0000;
	mel_filter_coefs[33][124] = 16'h0000;
	mel_filter_coefs[33][125] = 16'h0000;
	mel_filter_coefs[33][126] = 16'h0000;
	mel_filter_coefs[33][127] = 16'h0000;
	mel_filter_coefs[33][128] = 16'h0000;
	mel_filter_coefs[33][129] = 16'h0000;
	mel_filter_coefs[33][130] = 16'h0000;
	mel_filter_coefs[33][131] = 16'h0000;
	mel_filter_coefs[33][132] = 16'h0000;
	mel_filter_coefs[33][133] = 16'h0000;
	mel_filter_coefs[33][134] = 16'h0000;
	mel_filter_coefs[33][135] = 16'h0000;
	mel_filter_coefs[33][136] = 16'h0000;
	mel_filter_coefs[33][137] = 16'h0000;
	mel_filter_coefs[33][138] = 16'h0000;
	mel_filter_coefs[33][139] = 16'h0000;
	mel_filter_coefs[33][140] = 16'h0000;
	mel_filter_coefs[33][141] = 16'h0000;
	mel_filter_coefs[33][142] = 16'h0000;
	mel_filter_coefs[33][143] = 16'h0000;
	mel_filter_coefs[33][144] = 16'h0000;
	mel_filter_coefs[33][145] = 16'h0000;
	mel_filter_coefs[33][146] = 16'h0000;
	mel_filter_coefs[33][147] = 16'h0000;
	mel_filter_coefs[33][148] = 16'h087E;
	mel_filter_coefs[33][149] = 16'h1466;
	mel_filter_coefs[33][150] = 16'h204E;
	mel_filter_coefs[33][151] = 16'h2C36;
	mel_filter_coefs[33][152] = 16'h381D;
	mel_filter_coefs[33][153] = 16'h4405;
	mel_filter_coefs[33][154] = 16'h4FED;
	mel_filter_coefs[33][155] = 16'h5BD5;
	mel_filter_coefs[33][156] = 16'h67BD;
	mel_filter_coefs[33][157] = 16'h73A5;
	mel_filter_coefs[33][158] = 16'h7F8D;
	mel_filter_coefs[33][159] = 16'h753A;
	mel_filter_coefs[33][160] = 16'h6A08;
	mel_filter_coefs[33][161] = 16'h5ED6;
	mel_filter_coefs[33][162] = 16'h53A4;
	mel_filter_coefs[33][163] = 16'h4872;
	mel_filter_coefs[33][164] = 16'h3D40;
	mel_filter_coefs[33][165] = 16'h320D;
	mel_filter_coefs[33][166] = 16'h26DB;
	mel_filter_coefs[33][167] = 16'h1BA9;
	mel_filter_coefs[33][168] = 16'h1077;
	mel_filter_coefs[33][169] = 16'h0545;
	mel_filter_coefs[33][170] = 16'h0000;
	mel_filter_coefs[33][171] = 16'h0000;
	mel_filter_coefs[33][172] = 16'h0000;
	mel_filter_coefs[33][173] = 16'h0000;
	mel_filter_coefs[33][174] = 16'h0000;
	mel_filter_coefs[33][175] = 16'h0000;
	mel_filter_coefs[33][176] = 16'h0000;
	mel_filter_coefs[33][177] = 16'h0000;
	mel_filter_coefs[33][178] = 16'h0000;
	mel_filter_coefs[33][179] = 16'h0000;
	mel_filter_coefs[33][180] = 16'h0000;
	mel_filter_coefs[33][181] = 16'h0000;
	mel_filter_coefs[33][182] = 16'h0000;
	mel_filter_coefs[33][183] = 16'h0000;
	mel_filter_coefs[33][184] = 16'h0000;
	mel_filter_coefs[33][185] = 16'h0000;
	mel_filter_coefs[33][186] = 16'h0000;
	mel_filter_coefs[33][187] = 16'h0000;
	mel_filter_coefs[33][188] = 16'h0000;
	mel_filter_coefs[33][189] = 16'h0000;
	mel_filter_coefs[33][190] = 16'h0000;
	mel_filter_coefs[33][191] = 16'h0000;
	mel_filter_coefs[33][192] = 16'h0000;
	mel_filter_coefs[33][193] = 16'h0000;
	mel_filter_coefs[33][194] = 16'h0000;
	mel_filter_coefs[33][195] = 16'h0000;
	mel_filter_coefs[33][196] = 16'h0000;
	mel_filter_coefs[33][197] = 16'h0000;
	mel_filter_coefs[33][198] = 16'h0000;
	mel_filter_coefs[33][199] = 16'h0000;
	mel_filter_coefs[33][200] = 16'h0000;
	mel_filter_coefs[33][201] = 16'h0000;
	mel_filter_coefs[33][202] = 16'h0000;
	mel_filter_coefs[33][203] = 16'h0000;
	mel_filter_coefs[33][204] = 16'h0000;
	mel_filter_coefs[33][205] = 16'h0000;
	mel_filter_coefs[33][206] = 16'h0000;
	mel_filter_coefs[33][207] = 16'h0000;
	mel_filter_coefs[33][208] = 16'h0000;
	mel_filter_coefs[33][209] = 16'h0000;
	mel_filter_coefs[33][210] = 16'h0000;
	mel_filter_coefs[33][211] = 16'h0000;
	mel_filter_coefs[33][212] = 16'h0000;
	mel_filter_coefs[33][213] = 16'h0000;
	mel_filter_coefs[33][214] = 16'h0000;
	mel_filter_coefs[33][215] = 16'h0000;
	mel_filter_coefs[33][216] = 16'h0000;
	mel_filter_coefs[33][217] = 16'h0000;
	mel_filter_coefs[33][218] = 16'h0000;
	mel_filter_coefs[33][219] = 16'h0000;
	mel_filter_coefs[33][220] = 16'h0000;
	mel_filter_coefs[33][221] = 16'h0000;
	mel_filter_coefs[33][222] = 16'h0000;
	mel_filter_coefs[33][223] = 16'h0000;
	mel_filter_coefs[33][224] = 16'h0000;
	mel_filter_coefs[33][225] = 16'h0000;
	mel_filter_coefs[33][226] = 16'h0000;
	mel_filter_coefs[33][227] = 16'h0000;
	mel_filter_coefs[33][228] = 16'h0000;
	mel_filter_coefs[33][229] = 16'h0000;
	mel_filter_coefs[33][230] = 16'h0000;
	mel_filter_coefs[33][231] = 16'h0000;
	mel_filter_coefs[33][232] = 16'h0000;
	mel_filter_coefs[33][233] = 16'h0000;
	mel_filter_coefs[33][234] = 16'h0000;
	mel_filter_coefs[33][235] = 16'h0000;
	mel_filter_coefs[33][236] = 16'h0000;
	mel_filter_coefs[33][237] = 16'h0000;
	mel_filter_coefs[33][238] = 16'h0000;
	mel_filter_coefs[33][239] = 16'h0000;
	mel_filter_coefs[33][240] = 16'h0000;
	mel_filter_coefs[33][241] = 16'h0000;
	mel_filter_coefs[33][242] = 16'h0000;
	mel_filter_coefs[33][243] = 16'h0000;
	mel_filter_coefs[33][244] = 16'h0000;
	mel_filter_coefs[33][245] = 16'h0000;
	mel_filter_coefs[33][246] = 16'h0000;
	mel_filter_coefs[33][247] = 16'h0000;
	mel_filter_coefs[33][248] = 16'h0000;
	mel_filter_coefs[33][249] = 16'h0000;
	mel_filter_coefs[33][250] = 16'h0000;
	mel_filter_coefs[33][251] = 16'h0000;
	mel_filter_coefs[33][252] = 16'h0000;
	mel_filter_coefs[33][253] = 16'h0000;
	mel_filter_coefs[33][254] = 16'h0000;
	mel_filter_coefs[33][255] = 16'h0000;
	mel_filter_coefs[34][0] = 16'h0000;
	mel_filter_coefs[34][1] = 16'h0000;
	mel_filter_coefs[34][2] = 16'h0000;
	mel_filter_coefs[34][3] = 16'h0000;
	mel_filter_coefs[34][4] = 16'h0000;
	mel_filter_coefs[34][5] = 16'h0000;
	mel_filter_coefs[34][6] = 16'h0000;
	mel_filter_coefs[34][7] = 16'h0000;
	mel_filter_coefs[34][8] = 16'h0000;
	mel_filter_coefs[34][9] = 16'h0000;
	mel_filter_coefs[34][10] = 16'h0000;
	mel_filter_coefs[34][11] = 16'h0000;
	mel_filter_coefs[34][12] = 16'h0000;
	mel_filter_coefs[34][13] = 16'h0000;
	mel_filter_coefs[34][14] = 16'h0000;
	mel_filter_coefs[34][15] = 16'h0000;
	mel_filter_coefs[34][16] = 16'h0000;
	mel_filter_coefs[34][17] = 16'h0000;
	mel_filter_coefs[34][18] = 16'h0000;
	mel_filter_coefs[34][19] = 16'h0000;
	mel_filter_coefs[34][20] = 16'h0000;
	mel_filter_coefs[34][21] = 16'h0000;
	mel_filter_coefs[34][22] = 16'h0000;
	mel_filter_coefs[34][23] = 16'h0000;
	mel_filter_coefs[34][24] = 16'h0000;
	mel_filter_coefs[34][25] = 16'h0000;
	mel_filter_coefs[34][26] = 16'h0000;
	mel_filter_coefs[34][27] = 16'h0000;
	mel_filter_coefs[34][28] = 16'h0000;
	mel_filter_coefs[34][29] = 16'h0000;
	mel_filter_coefs[34][30] = 16'h0000;
	mel_filter_coefs[34][31] = 16'h0000;
	mel_filter_coefs[34][32] = 16'h0000;
	mel_filter_coefs[34][33] = 16'h0000;
	mel_filter_coefs[34][34] = 16'h0000;
	mel_filter_coefs[34][35] = 16'h0000;
	mel_filter_coefs[34][36] = 16'h0000;
	mel_filter_coefs[34][37] = 16'h0000;
	mel_filter_coefs[34][38] = 16'h0000;
	mel_filter_coefs[34][39] = 16'h0000;
	mel_filter_coefs[34][40] = 16'h0000;
	mel_filter_coefs[34][41] = 16'h0000;
	mel_filter_coefs[34][42] = 16'h0000;
	mel_filter_coefs[34][43] = 16'h0000;
	mel_filter_coefs[34][44] = 16'h0000;
	mel_filter_coefs[34][45] = 16'h0000;
	mel_filter_coefs[34][46] = 16'h0000;
	mel_filter_coefs[34][47] = 16'h0000;
	mel_filter_coefs[34][48] = 16'h0000;
	mel_filter_coefs[34][49] = 16'h0000;
	mel_filter_coefs[34][50] = 16'h0000;
	mel_filter_coefs[34][51] = 16'h0000;
	mel_filter_coefs[34][52] = 16'h0000;
	mel_filter_coefs[34][53] = 16'h0000;
	mel_filter_coefs[34][54] = 16'h0000;
	mel_filter_coefs[34][55] = 16'h0000;
	mel_filter_coefs[34][56] = 16'h0000;
	mel_filter_coefs[34][57] = 16'h0000;
	mel_filter_coefs[34][58] = 16'h0000;
	mel_filter_coefs[34][59] = 16'h0000;
	mel_filter_coefs[34][60] = 16'h0000;
	mel_filter_coefs[34][61] = 16'h0000;
	mel_filter_coefs[34][62] = 16'h0000;
	mel_filter_coefs[34][63] = 16'h0000;
	mel_filter_coefs[34][64] = 16'h0000;
	mel_filter_coefs[34][65] = 16'h0000;
	mel_filter_coefs[34][66] = 16'h0000;
	mel_filter_coefs[34][67] = 16'h0000;
	mel_filter_coefs[34][68] = 16'h0000;
	mel_filter_coefs[34][69] = 16'h0000;
	mel_filter_coefs[34][70] = 16'h0000;
	mel_filter_coefs[34][71] = 16'h0000;
	mel_filter_coefs[34][72] = 16'h0000;
	mel_filter_coefs[34][73] = 16'h0000;
	mel_filter_coefs[34][74] = 16'h0000;
	mel_filter_coefs[34][75] = 16'h0000;
	mel_filter_coefs[34][76] = 16'h0000;
	mel_filter_coefs[34][77] = 16'h0000;
	mel_filter_coefs[34][78] = 16'h0000;
	mel_filter_coefs[34][79] = 16'h0000;
	mel_filter_coefs[34][80] = 16'h0000;
	mel_filter_coefs[34][81] = 16'h0000;
	mel_filter_coefs[34][82] = 16'h0000;
	mel_filter_coefs[34][83] = 16'h0000;
	mel_filter_coefs[34][84] = 16'h0000;
	mel_filter_coefs[34][85] = 16'h0000;
	mel_filter_coefs[34][86] = 16'h0000;
	mel_filter_coefs[34][87] = 16'h0000;
	mel_filter_coefs[34][88] = 16'h0000;
	mel_filter_coefs[34][89] = 16'h0000;
	mel_filter_coefs[34][90] = 16'h0000;
	mel_filter_coefs[34][91] = 16'h0000;
	mel_filter_coefs[34][92] = 16'h0000;
	mel_filter_coefs[34][93] = 16'h0000;
	mel_filter_coefs[34][94] = 16'h0000;
	mel_filter_coefs[34][95] = 16'h0000;
	mel_filter_coefs[34][96] = 16'h0000;
	mel_filter_coefs[34][97] = 16'h0000;
	mel_filter_coefs[34][98] = 16'h0000;
	mel_filter_coefs[34][99] = 16'h0000;
	mel_filter_coefs[34][100] = 16'h0000;
	mel_filter_coefs[34][101] = 16'h0000;
	mel_filter_coefs[34][102] = 16'h0000;
	mel_filter_coefs[34][103] = 16'h0000;
	mel_filter_coefs[34][104] = 16'h0000;
	mel_filter_coefs[34][105] = 16'h0000;
	mel_filter_coefs[34][106] = 16'h0000;
	mel_filter_coefs[34][107] = 16'h0000;
	mel_filter_coefs[34][108] = 16'h0000;
	mel_filter_coefs[34][109] = 16'h0000;
	mel_filter_coefs[34][110] = 16'h0000;
	mel_filter_coefs[34][111] = 16'h0000;
	mel_filter_coefs[34][112] = 16'h0000;
	mel_filter_coefs[34][113] = 16'h0000;
	mel_filter_coefs[34][114] = 16'h0000;
	mel_filter_coefs[34][115] = 16'h0000;
	mel_filter_coefs[34][116] = 16'h0000;
	mel_filter_coefs[34][117] = 16'h0000;
	mel_filter_coefs[34][118] = 16'h0000;
	mel_filter_coefs[34][119] = 16'h0000;
	mel_filter_coefs[34][120] = 16'h0000;
	mel_filter_coefs[34][121] = 16'h0000;
	mel_filter_coefs[34][122] = 16'h0000;
	mel_filter_coefs[34][123] = 16'h0000;
	mel_filter_coefs[34][124] = 16'h0000;
	mel_filter_coefs[34][125] = 16'h0000;
	mel_filter_coefs[34][126] = 16'h0000;
	mel_filter_coefs[34][127] = 16'h0000;
	mel_filter_coefs[34][128] = 16'h0000;
	mel_filter_coefs[34][129] = 16'h0000;
	mel_filter_coefs[34][130] = 16'h0000;
	mel_filter_coefs[34][131] = 16'h0000;
	mel_filter_coefs[34][132] = 16'h0000;
	mel_filter_coefs[34][133] = 16'h0000;
	mel_filter_coefs[34][134] = 16'h0000;
	mel_filter_coefs[34][135] = 16'h0000;
	mel_filter_coefs[34][136] = 16'h0000;
	mel_filter_coefs[34][137] = 16'h0000;
	mel_filter_coefs[34][138] = 16'h0000;
	mel_filter_coefs[34][139] = 16'h0000;
	mel_filter_coefs[34][140] = 16'h0000;
	mel_filter_coefs[34][141] = 16'h0000;
	mel_filter_coefs[34][142] = 16'h0000;
	mel_filter_coefs[34][143] = 16'h0000;
	mel_filter_coefs[34][144] = 16'h0000;
	mel_filter_coefs[34][145] = 16'h0000;
	mel_filter_coefs[34][146] = 16'h0000;
	mel_filter_coefs[34][147] = 16'h0000;
	mel_filter_coefs[34][148] = 16'h0000;
	mel_filter_coefs[34][149] = 16'h0000;
	mel_filter_coefs[34][150] = 16'h0000;
	mel_filter_coefs[34][151] = 16'h0000;
	mel_filter_coefs[34][152] = 16'h0000;
	mel_filter_coefs[34][153] = 16'h0000;
	mel_filter_coefs[34][154] = 16'h0000;
	mel_filter_coefs[34][155] = 16'h0000;
	mel_filter_coefs[34][156] = 16'h0000;
	mel_filter_coefs[34][157] = 16'h0000;
	mel_filter_coefs[34][158] = 16'h0000;
	mel_filter_coefs[34][159] = 16'h0AC6;
	mel_filter_coefs[34][160] = 16'h15F8;
	mel_filter_coefs[34][161] = 16'h212A;
	mel_filter_coefs[34][162] = 16'h2C5C;
	mel_filter_coefs[34][163] = 16'h378E;
	mel_filter_coefs[34][164] = 16'h42C0;
	mel_filter_coefs[34][165] = 16'h4DF3;
	mel_filter_coefs[34][166] = 16'h5925;
	mel_filter_coefs[34][167] = 16'h6457;
	mel_filter_coefs[34][168] = 16'h6F89;
	mel_filter_coefs[34][169] = 16'h7ABB;
	mel_filter_coefs[34][170] = 16'h7A6D;
	mel_filter_coefs[34][171] = 16'h6FE6;
	mel_filter_coefs[34][172] = 16'h655E;
	mel_filter_coefs[34][173] = 16'h5AD7;
	mel_filter_coefs[34][174] = 16'h5050;
	mel_filter_coefs[34][175] = 16'h45C8;
	mel_filter_coefs[34][176] = 16'h3B41;
	mel_filter_coefs[34][177] = 16'h30BA;
	mel_filter_coefs[34][178] = 16'h2633;
	mel_filter_coefs[34][179] = 16'h1BAB;
	mel_filter_coefs[34][180] = 16'h1124;
	mel_filter_coefs[34][181] = 16'h069D;
	mel_filter_coefs[34][182] = 16'h0000;
	mel_filter_coefs[34][183] = 16'h0000;
	mel_filter_coefs[34][184] = 16'h0000;
	mel_filter_coefs[34][185] = 16'h0000;
	mel_filter_coefs[34][186] = 16'h0000;
	mel_filter_coefs[34][187] = 16'h0000;
	mel_filter_coefs[34][188] = 16'h0000;
	mel_filter_coefs[34][189] = 16'h0000;
	mel_filter_coefs[34][190] = 16'h0000;
	mel_filter_coefs[34][191] = 16'h0000;
	mel_filter_coefs[34][192] = 16'h0000;
	mel_filter_coefs[34][193] = 16'h0000;
	mel_filter_coefs[34][194] = 16'h0000;
	mel_filter_coefs[34][195] = 16'h0000;
	mel_filter_coefs[34][196] = 16'h0000;
	mel_filter_coefs[34][197] = 16'h0000;
	mel_filter_coefs[34][198] = 16'h0000;
	mel_filter_coefs[34][199] = 16'h0000;
	mel_filter_coefs[34][200] = 16'h0000;
	mel_filter_coefs[34][201] = 16'h0000;
	mel_filter_coefs[34][202] = 16'h0000;
	mel_filter_coefs[34][203] = 16'h0000;
	mel_filter_coefs[34][204] = 16'h0000;
	mel_filter_coefs[34][205] = 16'h0000;
	mel_filter_coefs[34][206] = 16'h0000;
	mel_filter_coefs[34][207] = 16'h0000;
	mel_filter_coefs[34][208] = 16'h0000;
	mel_filter_coefs[34][209] = 16'h0000;
	mel_filter_coefs[34][210] = 16'h0000;
	mel_filter_coefs[34][211] = 16'h0000;
	mel_filter_coefs[34][212] = 16'h0000;
	mel_filter_coefs[34][213] = 16'h0000;
	mel_filter_coefs[34][214] = 16'h0000;
	mel_filter_coefs[34][215] = 16'h0000;
	mel_filter_coefs[34][216] = 16'h0000;
	mel_filter_coefs[34][217] = 16'h0000;
	mel_filter_coefs[34][218] = 16'h0000;
	mel_filter_coefs[34][219] = 16'h0000;
	mel_filter_coefs[34][220] = 16'h0000;
	mel_filter_coefs[34][221] = 16'h0000;
	mel_filter_coefs[34][222] = 16'h0000;
	mel_filter_coefs[34][223] = 16'h0000;
	mel_filter_coefs[34][224] = 16'h0000;
	mel_filter_coefs[34][225] = 16'h0000;
	mel_filter_coefs[34][226] = 16'h0000;
	mel_filter_coefs[34][227] = 16'h0000;
	mel_filter_coefs[34][228] = 16'h0000;
	mel_filter_coefs[34][229] = 16'h0000;
	mel_filter_coefs[34][230] = 16'h0000;
	mel_filter_coefs[34][231] = 16'h0000;
	mel_filter_coefs[34][232] = 16'h0000;
	mel_filter_coefs[34][233] = 16'h0000;
	mel_filter_coefs[34][234] = 16'h0000;
	mel_filter_coefs[34][235] = 16'h0000;
	mel_filter_coefs[34][236] = 16'h0000;
	mel_filter_coefs[34][237] = 16'h0000;
	mel_filter_coefs[34][238] = 16'h0000;
	mel_filter_coefs[34][239] = 16'h0000;
	mel_filter_coefs[34][240] = 16'h0000;
	mel_filter_coefs[34][241] = 16'h0000;
	mel_filter_coefs[34][242] = 16'h0000;
	mel_filter_coefs[34][243] = 16'h0000;
	mel_filter_coefs[34][244] = 16'h0000;
	mel_filter_coefs[34][245] = 16'h0000;
	mel_filter_coefs[34][246] = 16'h0000;
	mel_filter_coefs[34][247] = 16'h0000;
	mel_filter_coefs[34][248] = 16'h0000;
	mel_filter_coefs[34][249] = 16'h0000;
	mel_filter_coefs[34][250] = 16'h0000;
	mel_filter_coefs[34][251] = 16'h0000;
	mel_filter_coefs[34][252] = 16'h0000;
	mel_filter_coefs[34][253] = 16'h0000;
	mel_filter_coefs[34][254] = 16'h0000;
	mel_filter_coefs[34][255] = 16'h0000;
	mel_filter_coefs[35][0] = 16'h0000;
	mel_filter_coefs[35][1] = 16'h0000;
	mel_filter_coefs[35][2] = 16'h0000;
	mel_filter_coefs[35][3] = 16'h0000;
	mel_filter_coefs[35][4] = 16'h0000;
	mel_filter_coefs[35][5] = 16'h0000;
	mel_filter_coefs[35][6] = 16'h0000;
	mel_filter_coefs[35][7] = 16'h0000;
	mel_filter_coefs[35][8] = 16'h0000;
	mel_filter_coefs[35][9] = 16'h0000;
	mel_filter_coefs[35][10] = 16'h0000;
	mel_filter_coefs[35][11] = 16'h0000;
	mel_filter_coefs[35][12] = 16'h0000;
	mel_filter_coefs[35][13] = 16'h0000;
	mel_filter_coefs[35][14] = 16'h0000;
	mel_filter_coefs[35][15] = 16'h0000;
	mel_filter_coefs[35][16] = 16'h0000;
	mel_filter_coefs[35][17] = 16'h0000;
	mel_filter_coefs[35][18] = 16'h0000;
	mel_filter_coefs[35][19] = 16'h0000;
	mel_filter_coefs[35][20] = 16'h0000;
	mel_filter_coefs[35][21] = 16'h0000;
	mel_filter_coefs[35][22] = 16'h0000;
	mel_filter_coefs[35][23] = 16'h0000;
	mel_filter_coefs[35][24] = 16'h0000;
	mel_filter_coefs[35][25] = 16'h0000;
	mel_filter_coefs[35][26] = 16'h0000;
	mel_filter_coefs[35][27] = 16'h0000;
	mel_filter_coefs[35][28] = 16'h0000;
	mel_filter_coefs[35][29] = 16'h0000;
	mel_filter_coefs[35][30] = 16'h0000;
	mel_filter_coefs[35][31] = 16'h0000;
	mel_filter_coefs[35][32] = 16'h0000;
	mel_filter_coefs[35][33] = 16'h0000;
	mel_filter_coefs[35][34] = 16'h0000;
	mel_filter_coefs[35][35] = 16'h0000;
	mel_filter_coefs[35][36] = 16'h0000;
	mel_filter_coefs[35][37] = 16'h0000;
	mel_filter_coefs[35][38] = 16'h0000;
	mel_filter_coefs[35][39] = 16'h0000;
	mel_filter_coefs[35][40] = 16'h0000;
	mel_filter_coefs[35][41] = 16'h0000;
	mel_filter_coefs[35][42] = 16'h0000;
	mel_filter_coefs[35][43] = 16'h0000;
	mel_filter_coefs[35][44] = 16'h0000;
	mel_filter_coefs[35][45] = 16'h0000;
	mel_filter_coefs[35][46] = 16'h0000;
	mel_filter_coefs[35][47] = 16'h0000;
	mel_filter_coefs[35][48] = 16'h0000;
	mel_filter_coefs[35][49] = 16'h0000;
	mel_filter_coefs[35][50] = 16'h0000;
	mel_filter_coefs[35][51] = 16'h0000;
	mel_filter_coefs[35][52] = 16'h0000;
	mel_filter_coefs[35][53] = 16'h0000;
	mel_filter_coefs[35][54] = 16'h0000;
	mel_filter_coefs[35][55] = 16'h0000;
	mel_filter_coefs[35][56] = 16'h0000;
	mel_filter_coefs[35][57] = 16'h0000;
	mel_filter_coefs[35][58] = 16'h0000;
	mel_filter_coefs[35][59] = 16'h0000;
	mel_filter_coefs[35][60] = 16'h0000;
	mel_filter_coefs[35][61] = 16'h0000;
	mel_filter_coefs[35][62] = 16'h0000;
	mel_filter_coefs[35][63] = 16'h0000;
	mel_filter_coefs[35][64] = 16'h0000;
	mel_filter_coefs[35][65] = 16'h0000;
	mel_filter_coefs[35][66] = 16'h0000;
	mel_filter_coefs[35][67] = 16'h0000;
	mel_filter_coefs[35][68] = 16'h0000;
	mel_filter_coefs[35][69] = 16'h0000;
	mel_filter_coefs[35][70] = 16'h0000;
	mel_filter_coefs[35][71] = 16'h0000;
	mel_filter_coefs[35][72] = 16'h0000;
	mel_filter_coefs[35][73] = 16'h0000;
	mel_filter_coefs[35][74] = 16'h0000;
	mel_filter_coefs[35][75] = 16'h0000;
	mel_filter_coefs[35][76] = 16'h0000;
	mel_filter_coefs[35][77] = 16'h0000;
	mel_filter_coefs[35][78] = 16'h0000;
	mel_filter_coefs[35][79] = 16'h0000;
	mel_filter_coefs[35][80] = 16'h0000;
	mel_filter_coefs[35][81] = 16'h0000;
	mel_filter_coefs[35][82] = 16'h0000;
	mel_filter_coefs[35][83] = 16'h0000;
	mel_filter_coefs[35][84] = 16'h0000;
	mel_filter_coefs[35][85] = 16'h0000;
	mel_filter_coefs[35][86] = 16'h0000;
	mel_filter_coefs[35][87] = 16'h0000;
	mel_filter_coefs[35][88] = 16'h0000;
	mel_filter_coefs[35][89] = 16'h0000;
	mel_filter_coefs[35][90] = 16'h0000;
	mel_filter_coefs[35][91] = 16'h0000;
	mel_filter_coefs[35][92] = 16'h0000;
	mel_filter_coefs[35][93] = 16'h0000;
	mel_filter_coefs[35][94] = 16'h0000;
	mel_filter_coefs[35][95] = 16'h0000;
	mel_filter_coefs[35][96] = 16'h0000;
	mel_filter_coefs[35][97] = 16'h0000;
	mel_filter_coefs[35][98] = 16'h0000;
	mel_filter_coefs[35][99] = 16'h0000;
	mel_filter_coefs[35][100] = 16'h0000;
	mel_filter_coefs[35][101] = 16'h0000;
	mel_filter_coefs[35][102] = 16'h0000;
	mel_filter_coefs[35][103] = 16'h0000;
	mel_filter_coefs[35][104] = 16'h0000;
	mel_filter_coefs[35][105] = 16'h0000;
	mel_filter_coefs[35][106] = 16'h0000;
	mel_filter_coefs[35][107] = 16'h0000;
	mel_filter_coefs[35][108] = 16'h0000;
	mel_filter_coefs[35][109] = 16'h0000;
	mel_filter_coefs[35][110] = 16'h0000;
	mel_filter_coefs[35][111] = 16'h0000;
	mel_filter_coefs[35][112] = 16'h0000;
	mel_filter_coefs[35][113] = 16'h0000;
	mel_filter_coefs[35][114] = 16'h0000;
	mel_filter_coefs[35][115] = 16'h0000;
	mel_filter_coefs[35][116] = 16'h0000;
	mel_filter_coefs[35][117] = 16'h0000;
	mel_filter_coefs[35][118] = 16'h0000;
	mel_filter_coefs[35][119] = 16'h0000;
	mel_filter_coefs[35][120] = 16'h0000;
	mel_filter_coefs[35][121] = 16'h0000;
	mel_filter_coefs[35][122] = 16'h0000;
	mel_filter_coefs[35][123] = 16'h0000;
	mel_filter_coefs[35][124] = 16'h0000;
	mel_filter_coefs[35][125] = 16'h0000;
	mel_filter_coefs[35][126] = 16'h0000;
	mel_filter_coefs[35][127] = 16'h0000;
	mel_filter_coefs[35][128] = 16'h0000;
	mel_filter_coefs[35][129] = 16'h0000;
	mel_filter_coefs[35][130] = 16'h0000;
	mel_filter_coefs[35][131] = 16'h0000;
	mel_filter_coefs[35][132] = 16'h0000;
	mel_filter_coefs[35][133] = 16'h0000;
	mel_filter_coefs[35][134] = 16'h0000;
	mel_filter_coefs[35][135] = 16'h0000;
	mel_filter_coefs[35][136] = 16'h0000;
	mel_filter_coefs[35][137] = 16'h0000;
	mel_filter_coefs[35][138] = 16'h0000;
	mel_filter_coefs[35][139] = 16'h0000;
	mel_filter_coefs[35][140] = 16'h0000;
	mel_filter_coefs[35][141] = 16'h0000;
	mel_filter_coefs[35][142] = 16'h0000;
	mel_filter_coefs[35][143] = 16'h0000;
	mel_filter_coefs[35][144] = 16'h0000;
	mel_filter_coefs[35][145] = 16'h0000;
	mel_filter_coefs[35][146] = 16'h0000;
	mel_filter_coefs[35][147] = 16'h0000;
	mel_filter_coefs[35][148] = 16'h0000;
	mel_filter_coefs[35][149] = 16'h0000;
	mel_filter_coefs[35][150] = 16'h0000;
	mel_filter_coefs[35][151] = 16'h0000;
	mel_filter_coefs[35][152] = 16'h0000;
	mel_filter_coefs[35][153] = 16'h0000;
	mel_filter_coefs[35][154] = 16'h0000;
	mel_filter_coefs[35][155] = 16'h0000;
	mel_filter_coefs[35][156] = 16'h0000;
	mel_filter_coefs[35][157] = 16'h0000;
	mel_filter_coefs[35][158] = 16'h0000;
	mel_filter_coefs[35][159] = 16'h0000;
	mel_filter_coefs[35][160] = 16'h0000;
	mel_filter_coefs[35][161] = 16'h0000;
	mel_filter_coefs[35][162] = 16'h0000;
	mel_filter_coefs[35][163] = 16'h0000;
	mel_filter_coefs[35][164] = 16'h0000;
	mel_filter_coefs[35][165] = 16'h0000;
	mel_filter_coefs[35][166] = 16'h0000;
	mel_filter_coefs[35][167] = 16'h0000;
	mel_filter_coefs[35][168] = 16'h0000;
	mel_filter_coefs[35][169] = 16'h0000;
	mel_filter_coefs[35][170] = 16'h0593;
	mel_filter_coefs[35][171] = 16'h101A;
	mel_filter_coefs[35][172] = 16'h1AA2;
	mel_filter_coefs[35][173] = 16'h2529;
	mel_filter_coefs[35][174] = 16'h2FB0;
	mel_filter_coefs[35][175] = 16'h3A38;
	mel_filter_coefs[35][176] = 16'h44BF;
	mel_filter_coefs[35][177] = 16'h4F46;
	mel_filter_coefs[35][178] = 16'h59CD;
	mel_filter_coefs[35][179] = 16'h6455;
	mel_filter_coefs[35][180] = 16'h6EDC;
	mel_filter_coefs[35][181] = 16'h7963;
	mel_filter_coefs[35][182] = 16'h7C51;
	mel_filter_coefs[35][183] = 16'h726A;
	mel_filter_coefs[35][184] = 16'h6884;
	mel_filter_coefs[35][185] = 16'h5E9D;
	mel_filter_coefs[35][186] = 16'h54B7;
	mel_filter_coefs[35][187] = 16'h4AD0;
	mel_filter_coefs[35][188] = 16'h40E9;
	mel_filter_coefs[35][189] = 16'h3703;
	mel_filter_coefs[35][190] = 16'h2D1C;
	mel_filter_coefs[35][191] = 16'h2335;
	mel_filter_coefs[35][192] = 16'h194F;
	mel_filter_coefs[35][193] = 16'h0F68;
	mel_filter_coefs[35][194] = 16'h0581;
	mel_filter_coefs[35][195] = 16'h0000;
	mel_filter_coefs[35][196] = 16'h0000;
	mel_filter_coefs[35][197] = 16'h0000;
	mel_filter_coefs[35][198] = 16'h0000;
	mel_filter_coefs[35][199] = 16'h0000;
	mel_filter_coefs[35][200] = 16'h0000;
	mel_filter_coefs[35][201] = 16'h0000;
	mel_filter_coefs[35][202] = 16'h0000;
	mel_filter_coefs[35][203] = 16'h0000;
	mel_filter_coefs[35][204] = 16'h0000;
	mel_filter_coefs[35][205] = 16'h0000;
	mel_filter_coefs[35][206] = 16'h0000;
	mel_filter_coefs[35][207] = 16'h0000;
	mel_filter_coefs[35][208] = 16'h0000;
	mel_filter_coefs[35][209] = 16'h0000;
	mel_filter_coefs[35][210] = 16'h0000;
	mel_filter_coefs[35][211] = 16'h0000;
	mel_filter_coefs[35][212] = 16'h0000;
	mel_filter_coefs[35][213] = 16'h0000;
	mel_filter_coefs[35][214] = 16'h0000;
	mel_filter_coefs[35][215] = 16'h0000;
	mel_filter_coefs[35][216] = 16'h0000;
	mel_filter_coefs[35][217] = 16'h0000;
	mel_filter_coefs[35][218] = 16'h0000;
	mel_filter_coefs[35][219] = 16'h0000;
	mel_filter_coefs[35][220] = 16'h0000;
	mel_filter_coefs[35][221] = 16'h0000;
	mel_filter_coefs[35][222] = 16'h0000;
	mel_filter_coefs[35][223] = 16'h0000;
	mel_filter_coefs[35][224] = 16'h0000;
	mel_filter_coefs[35][225] = 16'h0000;
	mel_filter_coefs[35][226] = 16'h0000;
	mel_filter_coefs[35][227] = 16'h0000;
	mel_filter_coefs[35][228] = 16'h0000;
	mel_filter_coefs[35][229] = 16'h0000;
	mel_filter_coefs[35][230] = 16'h0000;
	mel_filter_coefs[35][231] = 16'h0000;
	mel_filter_coefs[35][232] = 16'h0000;
	mel_filter_coefs[35][233] = 16'h0000;
	mel_filter_coefs[35][234] = 16'h0000;
	mel_filter_coefs[35][235] = 16'h0000;
	mel_filter_coefs[35][236] = 16'h0000;
	mel_filter_coefs[35][237] = 16'h0000;
	mel_filter_coefs[35][238] = 16'h0000;
	mel_filter_coefs[35][239] = 16'h0000;
	mel_filter_coefs[35][240] = 16'h0000;
	mel_filter_coefs[35][241] = 16'h0000;
	mel_filter_coefs[35][242] = 16'h0000;
	mel_filter_coefs[35][243] = 16'h0000;
	mel_filter_coefs[35][244] = 16'h0000;
	mel_filter_coefs[35][245] = 16'h0000;
	mel_filter_coefs[35][246] = 16'h0000;
	mel_filter_coefs[35][247] = 16'h0000;
	mel_filter_coefs[35][248] = 16'h0000;
	mel_filter_coefs[35][249] = 16'h0000;
	mel_filter_coefs[35][250] = 16'h0000;
	mel_filter_coefs[35][251] = 16'h0000;
	mel_filter_coefs[35][252] = 16'h0000;
	mel_filter_coefs[35][253] = 16'h0000;
	mel_filter_coefs[35][254] = 16'h0000;
	mel_filter_coefs[35][255] = 16'h0000;
	mel_filter_coefs[36][0] = 16'h0000;
	mel_filter_coefs[36][1] = 16'h0000;
	mel_filter_coefs[36][2] = 16'h0000;
	mel_filter_coefs[36][3] = 16'h0000;
	mel_filter_coefs[36][4] = 16'h0000;
	mel_filter_coefs[36][5] = 16'h0000;
	mel_filter_coefs[36][6] = 16'h0000;
	mel_filter_coefs[36][7] = 16'h0000;
	mel_filter_coefs[36][8] = 16'h0000;
	mel_filter_coefs[36][9] = 16'h0000;
	mel_filter_coefs[36][10] = 16'h0000;
	mel_filter_coefs[36][11] = 16'h0000;
	mel_filter_coefs[36][12] = 16'h0000;
	mel_filter_coefs[36][13] = 16'h0000;
	mel_filter_coefs[36][14] = 16'h0000;
	mel_filter_coefs[36][15] = 16'h0000;
	mel_filter_coefs[36][16] = 16'h0000;
	mel_filter_coefs[36][17] = 16'h0000;
	mel_filter_coefs[36][18] = 16'h0000;
	mel_filter_coefs[36][19] = 16'h0000;
	mel_filter_coefs[36][20] = 16'h0000;
	mel_filter_coefs[36][21] = 16'h0000;
	mel_filter_coefs[36][22] = 16'h0000;
	mel_filter_coefs[36][23] = 16'h0000;
	mel_filter_coefs[36][24] = 16'h0000;
	mel_filter_coefs[36][25] = 16'h0000;
	mel_filter_coefs[36][26] = 16'h0000;
	mel_filter_coefs[36][27] = 16'h0000;
	mel_filter_coefs[36][28] = 16'h0000;
	mel_filter_coefs[36][29] = 16'h0000;
	mel_filter_coefs[36][30] = 16'h0000;
	mel_filter_coefs[36][31] = 16'h0000;
	mel_filter_coefs[36][32] = 16'h0000;
	mel_filter_coefs[36][33] = 16'h0000;
	mel_filter_coefs[36][34] = 16'h0000;
	mel_filter_coefs[36][35] = 16'h0000;
	mel_filter_coefs[36][36] = 16'h0000;
	mel_filter_coefs[36][37] = 16'h0000;
	mel_filter_coefs[36][38] = 16'h0000;
	mel_filter_coefs[36][39] = 16'h0000;
	mel_filter_coefs[36][40] = 16'h0000;
	mel_filter_coefs[36][41] = 16'h0000;
	mel_filter_coefs[36][42] = 16'h0000;
	mel_filter_coefs[36][43] = 16'h0000;
	mel_filter_coefs[36][44] = 16'h0000;
	mel_filter_coefs[36][45] = 16'h0000;
	mel_filter_coefs[36][46] = 16'h0000;
	mel_filter_coefs[36][47] = 16'h0000;
	mel_filter_coefs[36][48] = 16'h0000;
	mel_filter_coefs[36][49] = 16'h0000;
	mel_filter_coefs[36][50] = 16'h0000;
	mel_filter_coefs[36][51] = 16'h0000;
	mel_filter_coefs[36][52] = 16'h0000;
	mel_filter_coefs[36][53] = 16'h0000;
	mel_filter_coefs[36][54] = 16'h0000;
	mel_filter_coefs[36][55] = 16'h0000;
	mel_filter_coefs[36][56] = 16'h0000;
	mel_filter_coefs[36][57] = 16'h0000;
	mel_filter_coefs[36][58] = 16'h0000;
	mel_filter_coefs[36][59] = 16'h0000;
	mel_filter_coefs[36][60] = 16'h0000;
	mel_filter_coefs[36][61] = 16'h0000;
	mel_filter_coefs[36][62] = 16'h0000;
	mel_filter_coefs[36][63] = 16'h0000;
	mel_filter_coefs[36][64] = 16'h0000;
	mel_filter_coefs[36][65] = 16'h0000;
	mel_filter_coefs[36][66] = 16'h0000;
	mel_filter_coefs[36][67] = 16'h0000;
	mel_filter_coefs[36][68] = 16'h0000;
	mel_filter_coefs[36][69] = 16'h0000;
	mel_filter_coefs[36][70] = 16'h0000;
	mel_filter_coefs[36][71] = 16'h0000;
	mel_filter_coefs[36][72] = 16'h0000;
	mel_filter_coefs[36][73] = 16'h0000;
	mel_filter_coefs[36][74] = 16'h0000;
	mel_filter_coefs[36][75] = 16'h0000;
	mel_filter_coefs[36][76] = 16'h0000;
	mel_filter_coefs[36][77] = 16'h0000;
	mel_filter_coefs[36][78] = 16'h0000;
	mel_filter_coefs[36][79] = 16'h0000;
	mel_filter_coefs[36][80] = 16'h0000;
	mel_filter_coefs[36][81] = 16'h0000;
	mel_filter_coefs[36][82] = 16'h0000;
	mel_filter_coefs[36][83] = 16'h0000;
	mel_filter_coefs[36][84] = 16'h0000;
	mel_filter_coefs[36][85] = 16'h0000;
	mel_filter_coefs[36][86] = 16'h0000;
	mel_filter_coefs[36][87] = 16'h0000;
	mel_filter_coefs[36][88] = 16'h0000;
	mel_filter_coefs[36][89] = 16'h0000;
	mel_filter_coefs[36][90] = 16'h0000;
	mel_filter_coefs[36][91] = 16'h0000;
	mel_filter_coefs[36][92] = 16'h0000;
	mel_filter_coefs[36][93] = 16'h0000;
	mel_filter_coefs[36][94] = 16'h0000;
	mel_filter_coefs[36][95] = 16'h0000;
	mel_filter_coefs[36][96] = 16'h0000;
	mel_filter_coefs[36][97] = 16'h0000;
	mel_filter_coefs[36][98] = 16'h0000;
	mel_filter_coefs[36][99] = 16'h0000;
	mel_filter_coefs[36][100] = 16'h0000;
	mel_filter_coefs[36][101] = 16'h0000;
	mel_filter_coefs[36][102] = 16'h0000;
	mel_filter_coefs[36][103] = 16'h0000;
	mel_filter_coefs[36][104] = 16'h0000;
	mel_filter_coefs[36][105] = 16'h0000;
	mel_filter_coefs[36][106] = 16'h0000;
	mel_filter_coefs[36][107] = 16'h0000;
	mel_filter_coefs[36][108] = 16'h0000;
	mel_filter_coefs[36][109] = 16'h0000;
	mel_filter_coefs[36][110] = 16'h0000;
	mel_filter_coefs[36][111] = 16'h0000;
	mel_filter_coefs[36][112] = 16'h0000;
	mel_filter_coefs[36][113] = 16'h0000;
	mel_filter_coefs[36][114] = 16'h0000;
	mel_filter_coefs[36][115] = 16'h0000;
	mel_filter_coefs[36][116] = 16'h0000;
	mel_filter_coefs[36][117] = 16'h0000;
	mel_filter_coefs[36][118] = 16'h0000;
	mel_filter_coefs[36][119] = 16'h0000;
	mel_filter_coefs[36][120] = 16'h0000;
	mel_filter_coefs[36][121] = 16'h0000;
	mel_filter_coefs[36][122] = 16'h0000;
	mel_filter_coefs[36][123] = 16'h0000;
	mel_filter_coefs[36][124] = 16'h0000;
	mel_filter_coefs[36][125] = 16'h0000;
	mel_filter_coefs[36][126] = 16'h0000;
	mel_filter_coefs[36][127] = 16'h0000;
	mel_filter_coefs[36][128] = 16'h0000;
	mel_filter_coefs[36][129] = 16'h0000;
	mel_filter_coefs[36][130] = 16'h0000;
	mel_filter_coefs[36][131] = 16'h0000;
	mel_filter_coefs[36][132] = 16'h0000;
	mel_filter_coefs[36][133] = 16'h0000;
	mel_filter_coefs[36][134] = 16'h0000;
	mel_filter_coefs[36][135] = 16'h0000;
	mel_filter_coefs[36][136] = 16'h0000;
	mel_filter_coefs[36][137] = 16'h0000;
	mel_filter_coefs[36][138] = 16'h0000;
	mel_filter_coefs[36][139] = 16'h0000;
	mel_filter_coefs[36][140] = 16'h0000;
	mel_filter_coefs[36][141] = 16'h0000;
	mel_filter_coefs[36][142] = 16'h0000;
	mel_filter_coefs[36][143] = 16'h0000;
	mel_filter_coefs[36][144] = 16'h0000;
	mel_filter_coefs[36][145] = 16'h0000;
	mel_filter_coefs[36][146] = 16'h0000;
	mel_filter_coefs[36][147] = 16'h0000;
	mel_filter_coefs[36][148] = 16'h0000;
	mel_filter_coefs[36][149] = 16'h0000;
	mel_filter_coefs[36][150] = 16'h0000;
	mel_filter_coefs[36][151] = 16'h0000;
	mel_filter_coefs[36][152] = 16'h0000;
	mel_filter_coefs[36][153] = 16'h0000;
	mel_filter_coefs[36][154] = 16'h0000;
	mel_filter_coefs[36][155] = 16'h0000;
	mel_filter_coefs[36][156] = 16'h0000;
	mel_filter_coefs[36][157] = 16'h0000;
	mel_filter_coefs[36][158] = 16'h0000;
	mel_filter_coefs[36][159] = 16'h0000;
	mel_filter_coefs[36][160] = 16'h0000;
	mel_filter_coefs[36][161] = 16'h0000;
	mel_filter_coefs[36][162] = 16'h0000;
	mel_filter_coefs[36][163] = 16'h0000;
	mel_filter_coefs[36][164] = 16'h0000;
	mel_filter_coefs[36][165] = 16'h0000;
	mel_filter_coefs[36][166] = 16'h0000;
	mel_filter_coefs[36][167] = 16'h0000;
	mel_filter_coefs[36][168] = 16'h0000;
	mel_filter_coefs[36][169] = 16'h0000;
	mel_filter_coefs[36][170] = 16'h0000;
	mel_filter_coefs[36][171] = 16'h0000;
	mel_filter_coefs[36][172] = 16'h0000;
	mel_filter_coefs[36][173] = 16'h0000;
	mel_filter_coefs[36][174] = 16'h0000;
	mel_filter_coefs[36][175] = 16'h0000;
	mel_filter_coefs[36][176] = 16'h0000;
	mel_filter_coefs[36][177] = 16'h0000;
	mel_filter_coefs[36][178] = 16'h0000;
	mel_filter_coefs[36][179] = 16'h0000;
	mel_filter_coefs[36][180] = 16'h0000;
	mel_filter_coefs[36][181] = 16'h0000;
	mel_filter_coefs[36][182] = 16'h03AF;
	mel_filter_coefs[36][183] = 16'h0D96;
	mel_filter_coefs[36][184] = 16'h177C;
	mel_filter_coefs[36][185] = 16'h2163;
	mel_filter_coefs[36][186] = 16'h2B49;
	mel_filter_coefs[36][187] = 16'h3530;
	mel_filter_coefs[36][188] = 16'h3F17;
	mel_filter_coefs[36][189] = 16'h48FD;
	mel_filter_coefs[36][190] = 16'h52E4;
	mel_filter_coefs[36][191] = 16'h5CCB;
	mel_filter_coefs[36][192] = 16'h66B1;
	mel_filter_coefs[36][193] = 16'h7098;
	mel_filter_coefs[36][194] = 16'h7A7F;
	mel_filter_coefs[36][195] = 16'h7BDE;
	mel_filter_coefs[36][196] = 16'h728E;
	mel_filter_coefs[36][197] = 16'h693F;
	mel_filter_coefs[36][198] = 16'h5FEF;
	mel_filter_coefs[36][199] = 16'h56A0;
	mel_filter_coefs[36][200] = 16'h4D50;
	mel_filter_coefs[36][201] = 16'h4401;
	mel_filter_coefs[36][202] = 16'h3AB1;
	mel_filter_coefs[36][203] = 16'h3162;
	mel_filter_coefs[36][204] = 16'h2812;
	mel_filter_coefs[36][205] = 16'h1EC3;
	mel_filter_coefs[36][206] = 16'h1573;
	mel_filter_coefs[36][207] = 16'h0C23;
	mel_filter_coefs[36][208] = 16'h02D4;
	mel_filter_coefs[36][209] = 16'h0000;
	mel_filter_coefs[36][210] = 16'h0000;
	mel_filter_coefs[36][211] = 16'h0000;
	mel_filter_coefs[36][212] = 16'h0000;
	mel_filter_coefs[36][213] = 16'h0000;
	mel_filter_coefs[36][214] = 16'h0000;
	mel_filter_coefs[36][215] = 16'h0000;
	mel_filter_coefs[36][216] = 16'h0000;
	mel_filter_coefs[36][217] = 16'h0000;
	mel_filter_coefs[36][218] = 16'h0000;
	mel_filter_coefs[36][219] = 16'h0000;
	mel_filter_coefs[36][220] = 16'h0000;
	mel_filter_coefs[36][221] = 16'h0000;
	mel_filter_coefs[36][222] = 16'h0000;
	mel_filter_coefs[36][223] = 16'h0000;
	mel_filter_coefs[36][224] = 16'h0000;
	mel_filter_coefs[36][225] = 16'h0000;
	mel_filter_coefs[36][226] = 16'h0000;
	mel_filter_coefs[36][227] = 16'h0000;
	mel_filter_coefs[36][228] = 16'h0000;
	mel_filter_coefs[36][229] = 16'h0000;
	mel_filter_coefs[36][230] = 16'h0000;
	mel_filter_coefs[36][231] = 16'h0000;
	mel_filter_coefs[36][232] = 16'h0000;
	mel_filter_coefs[36][233] = 16'h0000;
	mel_filter_coefs[36][234] = 16'h0000;
	mel_filter_coefs[36][235] = 16'h0000;
	mel_filter_coefs[36][236] = 16'h0000;
	mel_filter_coefs[36][237] = 16'h0000;
	mel_filter_coefs[36][238] = 16'h0000;
	mel_filter_coefs[36][239] = 16'h0000;
	mel_filter_coefs[36][240] = 16'h0000;
	mel_filter_coefs[36][241] = 16'h0000;
	mel_filter_coefs[36][242] = 16'h0000;
	mel_filter_coefs[36][243] = 16'h0000;
	mel_filter_coefs[36][244] = 16'h0000;
	mel_filter_coefs[36][245] = 16'h0000;
	mel_filter_coefs[36][246] = 16'h0000;
	mel_filter_coefs[36][247] = 16'h0000;
	mel_filter_coefs[36][248] = 16'h0000;
	mel_filter_coefs[36][249] = 16'h0000;
	mel_filter_coefs[36][250] = 16'h0000;
	mel_filter_coefs[36][251] = 16'h0000;
	mel_filter_coefs[36][252] = 16'h0000;
	mel_filter_coefs[36][253] = 16'h0000;
	mel_filter_coefs[36][254] = 16'h0000;
	mel_filter_coefs[36][255] = 16'h0000;
	mel_filter_coefs[37][0] = 16'h0000;
	mel_filter_coefs[37][1] = 16'h0000;
	mel_filter_coefs[37][2] = 16'h0000;
	mel_filter_coefs[37][3] = 16'h0000;
	mel_filter_coefs[37][4] = 16'h0000;
	mel_filter_coefs[37][5] = 16'h0000;
	mel_filter_coefs[37][6] = 16'h0000;
	mel_filter_coefs[37][7] = 16'h0000;
	mel_filter_coefs[37][8] = 16'h0000;
	mel_filter_coefs[37][9] = 16'h0000;
	mel_filter_coefs[37][10] = 16'h0000;
	mel_filter_coefs[37][11] = 16'h0000;
	mel_filter_coefs[37][12] = 16'h0000;
	mel_filter_coefs[37][13] = 16'h0000;
	mel_filter_coefs[37][14] = 16'h0000;
	mel_filter_coefs[37][15] = 16'h0000;
	mel_filter_coefs[37][16] = 16'h0000;
	mel_filter_coefs[37][17] = 16'h0000;
	mel_filter_coefs[37][18] = 16'h0000;
	mel_filter_coefs[37][19] = 16'h0000;
	mel_filter_coefs[37][20] = 16'h0000;
	mel_filter_coefs[37][21] = 16'h0000;
	mel_filter_coefs[37][22] = 16'h0000;
	mel_filter_coefs[37][23] = 16'h0000;
	mel_filter_coefs[37][24] = 16'h0000;
	mel_filter_coefs[37][25] = 16'h0000;
	mel_filter_coefs[37][26] = 16'h0000;
	mel_filter_coefs[37][27] = 16'h0000;
	mel_filter_coefs[37][28] = 16'h0000;
	mel_filter_coefs[37][29] = 16'h0000;
	mel_filter_coefs[37][30] = 16'h0000;
	mel_filter_coefs[37][31] = 16'h0000;
	mel_filter_coefs[37][32] = 16'h0000;
	mel_filter_coefs[37][33] = 16'h0000;
	mel_filter_coefs[37][34] = 16'h0000;
	mel_filter_coefs[37][35] = 16'h0000;
	mel_filter_coefs[37][36] = 16'h0000;
	mel_filter_coefs[37][37] = 16'h0000;
	mel_filter_coefs[37][38] = 16'h0000;
	mel_filter_coefs[37][39] = 16'h0000;
	mel_filter_coefs[37][40] = 16'h0000;
	mel_filter_coefs[37][41] = 16'h0000;
	mel_filter_coefs[37][42] = 16'h0000;
	mel_filter_coefs[37][43] = 16'h0000;
	mel_filter_coefs[37][44] = 16'h0000;
	mel_filter_coefs[37][45] = 16'h0000;
	mel_filter_coefs[37][46] = 16'h0000;
	mel_filter_coefs[37][47] = 16'h0000;
	mel_filter_coefs[37][48] = 16'h0000;
	mel_filter_coefs[37][49] = 16'h0000;
	mel_filter_coefs[37][50] = 16'h0000;
	mel_filter_coefs[37][51] = 16'h0000;
	mel_filter_coefs[37][52] = 16'h0000;
	mel_filter_coefs[37][53] = 16'h0000;
	mel_filter_coefs[37][54] = 16'h0000;
	mel_filter_coefs[37][55] = 16'h0000;
	mel_filter_coefs[37][56] = 16'h0000;
	mel_filter_coefs[37][57] = 16'h0000;
	mel_filter_coefs[37][58] = 16'h0000;
	mel_filter_coefs[37][59] = 16'h0000;
	mel_filter_coefs[37][60] = 16'h0000;
	mel_filter_coefs[37][61] = 16'h0000;
	mel_filter_coefs[37][62] = 16'h0000;
	mel_filter_coefs[37][63] = 16'h0000;
	mel_filter_coefs[37][64] = 16'h0000;
	mel_filter_coefs[37][65] = 16'h0000;
	mel_filter_coefs[37][66] = 16'h0000;
	mel_filter_coefs[37][67] = 16'h0000;
	mel_filter_coefs[37][68] = 16'h0000;
	mel_filter_coefs[37][69] = 16'h0000;
	mel_filter_coefs[37][70] = 16'h0000;
	mel_filter_coefs[37][71] = 16'h0000;
	mel_filter_coefs[37][72] = 16'h0000;
	mel_filter_coefs[37][73] = 16'h0000;
	mel_filter_coefs[37][74] = 16'h0000;
	mel_filter_coefs[37][75] = 16'h0000;
	mel_filter_coefs[37][76] = 16'h0000;
	mel_filter_coefs[37][77] = 16'h0000;
	mel_filter_coefs[37][78] = 16'h0000;
	mel_filter_coefs[37][79] = 16'h0000;
	mel_filter_coefs[37][80] = 16'h0000;
	mel_filter_coefs[37][81] = 16'h0000;
	mel_filter_coefs[37][82] = 16'h0000;
	mel_filter_coefs[37][83] = 16'h0000;
	mel_filter_coefs[37][84] = 16'h0000;
	mel_filter_coefs[37][85] = 16'h0000;
	mel_filter_coefs[37][86] = 16'h0000;
	mel_filter_coefs[37][87] = 16'h0000;
	mel_filter_coefs[37][88] = 16'h0000;
	mel_filter_coefs[37][89] = 16'h0000;
	mel_filter_coefs[37][90] = 16'h0000;
	mel_filter_coefs[37][91] = 16'h0000;
	mel_filter_coefs[37][92] = 16'h0000;
	mel_filter_coefs[37][93] = 16'h0000;
	mel_filter_coefs[37][94] = 16'h0000;
	mel_filter_coefs[37][95] = 16'h0000;
	mel_filter_coefs[37][96] = 16'h0000;
	mel_filter_coefs[37][97] = 16'h0000;
	mel_filter_coefs[37][98] = 16'h0000;
	mel_filter_coefs[37][99] = 16'h0000;
	mel_filter_coefs[37][100] = 16'h0000;
	mel_filter_coefs[37][101] = 16'h0000;
	mel_filter_coefs[37][102] = 16'h0000;
	mel_filter_coefs[37][103] = 16'h0000;
	mel_filter_coefs[37][104] = 16'h0000;
	mel_filter_coefs[37][105] = 16'h0000;
	mel_filter_coefs[37][106] = 16'h0000;
	mel_filter_coefs[37][107] = 16'h0000;
	mel_filter_coefs[37][108] = 16'h0000;
	mel_filter_coefs[37][109] = 16'h0000;
	mel_filter_coefs[37][110] = 16'h0000;
	mel_filter_coefs[37][111] = 16'h0000;
	mel_filter_coefs[37][112] = 16'h0000;
	mel_filter_coefs[37][113] = 16'h0000;
	mel_filter_coefs[37][114] = 16'h0000;
	mel_filter_coefs[37][115] = 16'h0000;
	mel_filter_coefs[37][116] = 16'h0000;
	mel_filter_coefs[37][117] = 16'h0000;
	mel_filter_coefs[37][118] = 16'h0000;
	mel_filter_coefs[37][119] = 16'h0000;
	mel_filter_coefs[37][120] = 16'h0000;
	mel_filter_coefs[37][121] = 16'h0000;
	mel_filter_coefs[37][122] = 16'h0000;
	mel_filter_coefs[37][123] = 16'h0000;
	mel_filter_coefs[37][124] = 16'h0000;
	mel_filter_coefs[37][125] = 16'h0000;
	mel_filter_coefs[37][126] = 16'h0000;
	mel_filter_coefs[37][127] = 16'h0000;
	mel_filter_coefs[37][128] = 16'h0000;
	mel_filter_coefs[37][129] = 16'h0000;
	mel_filter_coefs[37][130] = 16'h0000;
	mel_filter_coefs[37][131] = 16'h0000;
	mel_filter_coefs[37][132] = 16'h0000;
	mel_filter_coefs[37][133] = 16'h0000;
	mel_filter_coefs[37][134] = 16'h0000;
	mel_filter_coefs[37][135] = 16'h0000;
	mel_filter_coefs[37][136] = 16'h0000;
	mel_filter_coefs[37][137] = 16'h0000;
	mel_filter_coefs[37][138] = 16'h0000;
	mel_filter_coefs[37][139] = 16'h0000;
	mel_filter_coefs[37][140] = 16'h0000;
	mel_filter_coefs[37][141] = 16'h0000;
	mel_filter_coefs[37][142] = 16'h0000;
	mel_filter_coefs[37][143] = 16'h0000;
	mel_filter_coefs[37][144] = 16'h0000;
	mel_filter_coefs[37][145] = 16'h0000;
	mel_filter_coefs[37][146] = 16'h0000;
	mel_filter_coefs[37][147] = 16'h0000;
	mel_filter_coefs[37][148] = 16'h0000;
	mel_filter_coefs[37][149] = 16'h0000;
	mel_filter_coefs[37][150] = 16'h0000;
	mel_filter_coefs[37][151] = 16'h0000;
	mel_filter_coefs[37][152] = 16'h0000;
	mel_filter_coefs[37][153] = 16'h0000;
	mel_filter_coefs[37][154] = 16'h0000;
	mel_filter_coefs[37][155] = 16'h0000;
	mel_filter_coefs[37][156] = 16'h0000;
	mel_filter_coefs[37][157] = 16'h0000;
	mel_filter_coefs[37][158] = 16'h0000;
	mel_filter_coefs[37][159] = 16'h0000;
	mel_filter_coefs[37][160] = 16'h0000;
	mel_filter_coefs[37][161] = 16'h0000;
	mel_filter_coefs[37][162] = 16'h0000;
	mel_filter_coefs[37][163] = 16'h0000;
	mel_filter_coefs[37][164] = 16'h0000;
	mel_filter_coefs[37][165] = 16'h0000;
	mel_filter_coefs[37][166] = 16'h0000;
	mel_filter_coefs[37][167] = 16'h0000;
	mel_filter_coefs[37][168] = 16'h0000;
	mel_filter_coefs[37][169] = 16'h0000;
	mel_filter_coefs[37][170] = 16'h0000;
	mel_filter_coefs[37][171] = 16'h0000;
	mel_filter_coefs[37][172] = 16'h0000;
	mel_filter_coefs[37][173] = 16'h0000;
	mel_filter_coefs[37][174] = 16'h0000;
	mel_filter_coefs[37][175] = 16'h0000;
	mel_filter_coefs[37][176] = 16'h0000;
	mel_filter_coefs[37][177] = 16'h0000;
	mel_filter_coefs[37][178] = 16'h0000;
	mel_filter_coefs[37][179] = 16'h0000;
	mel_filter_coefs[37][180] = 16'h0000;
	mel_filter_coefs[37][181] = 16'h0000;
	mel_filter_coefs[37][182] = 16'h0000;
	mel_filter_coefs[37][183] = 16'h0000;
	mel_filter_coefs[37][184] = 16'h0000;
	mel_filter_coefs[37][185] = 16'h0000;
	mel_filter_coefs[37][186] = 16'h0000;
	mel_filter_coefs[37][187] = 16'h0000;
	mel_filter_coefs[37][188] = 16'h0000;
	mel_filter_coefs[37][189] = 16'h0000;
	mel_filter_coefs[37][190] = 16'h0000;
	mel_filter_coefs[37][191] = 16'h0000;
	mel_filter_coefs[37][192] = 16'h0000;
	mel_filter_coefs[37][193] = 16'h0000;
	mel_filter_coefs[37][194] = 16'h0000;
	mel_filter_coefs[37][195] = 16'h0422;
	mel_filter_coefs[37][196] = 16'h0D72;
	mel_filter_coefs[37][197] = 16'h16C1;
	mel_filter_coefs[37][198] = 16'h2011;
	mel_filter_coefs[37][199] = 16'h2960;
	mel_filter_coefs[37][200] = 16'h32B0;
	mel_filter_coefs[37][201] = 16'h3BFF;
	mel_filter_coefs[37][202] = 16'h454F;
	mel_filter_coefs[37][203] = 16'h4E9E;
	mel_filter_coefs[37][204] = 16'h57EE;
	mel_filter_coefs[37][205] = 16'h613D;
	mel_filter_coefs[37][206] = 16'h6A8D;
	mel_filter_coefs[37][207] = 16'h73DD;
	mel_filter_coefs[37][208] = 16'h7D2C;
	mel_filter_coefs[37][209] = 16'h79E7;
	mel_filter_coefs[37][210] = 16'h7126;
	mel_filter_coefs[37][211] = 16'h6864;
	mel_filter_coefs[37][212] = 16'h5FA3;
	mel_filter_coefs[37][213] = 16'h56E2;
	mel_filter_coefs[37][214] = 16'h4E20;
	mel_filter_coefs[37][215] = 16'h455F;
	mel_filter_coefs[37][216] = 16'h3C9D;
	mel_filter_coefs[37][217] = 16'h33DC;
	mel_filter_coefs[37][218] = 16'h2B1A;
	mel_filter_coefs[37][219] = 16'h2259;
	mel_filter_coefs[37][220] = 16'h1997;
	mel_filter_coefs[37][221] = 16'h10D6;
	mel_filter_coefs[37][222] = 16'h0814;
	mel_filter_coefs[37][223] = 16'h0000;
	mel_filter_coefs[37][224] = 16'h0000;
	mel_filter_coefs[37][225] = 16'h0000;
	mel_filter_coefs[37][226] = 16'h0000;
	mel_filter_coefs[37][227] = 16'h0000;
	mel_filter_coefs[37][228] = 16'h0000;
	mel_filter_coefs[37][229] = 16'h0000;
	mel_filter_coefs[37][230] = 16'h0000;
	mel_filter_coefs[37][231] = 16'h0000;
	mel_filter_coefs[37][232] = 16'h0000;
	mel_filter_coefs[37][233] = 16'h0000;
	mel_filter_coefs[37][234] = 16'h0000;
	mel_filter_coefs[37][235] = 16'h0000;
	mel_filter_coefs[37][236] = 16'h0000;
	mel_filter_coefs[37][237] = 16'h0000;
	mel_filter_coefs[37][238] = 16'h0000;
	mel_filter_coefs[37][239] = 16'h0000;
	mel_filter_coefs[37][240] = 16'h0000;
	mel_filter_coefs[37][241] = 16'h0000;
	mel_filter_coefs[37][242] = 16'h0000;
	mel_filter_coefs[37][243] = 16'h0000;
	mel_filter_coefs[37][244] = 16'h0000;
	mel_filter_coefs[37][245] = 16'h0000;
	mel_filter_coefs[37][246] = 16'h0000;
	mel_filter_coefs[37][247] = 16'h0000;
	mel_filter_coefs[37][248] = 16'h0000;
	mel_filter_coefs[37][249] = 16'h0000;
	mel_filter_coefs[37][250] = 16'h0000;
	mel_filter_coefs[37][251] = 16'h0000;
	mel_filter_coefs[37][252] = 16'h0000;
	mel_filter_coefs[37][253] = 16'h0000;
	mel_filter_coefs[37][254] = 16'h0000;
	mel_filter_coefs[37][255] = 16'h0000;
	mel_filter_coefs[38][0] = 16'h0000;
	mel_filter_coefs[38][1] = 16'h0000;
	mel_filter_coefs[38][2] = 16'h0000;
	mel_filter_coefs[38][3] = 16'h0000;
	mel_filter_coefs[38][4] = 16'h0000;
	mel_filter_coefs[38][5] = 16'h0000;
	mel_filter_coefs[38][6] = 16'h0000;
	mel_filter_coefs[38][7] = 16'h0000;
	mel_filter_coefs[38][8] = 16'h0000;
	mel_filter_coefs[38][9] = 16'h0000;
	mel_filter_coefs[38][10] = 16'h0000;
	mel_filter_coefs[38][11] = 16'h0000;
	mel_filter_coefs[38][12] = 16'h0000;
	mel_filter_coefs[38][13] = 16'h0000;
	mel_filter_coefs[38][14] = 16'h0000;
	mel_filter_coefs[38][15] = 16'h0000;
	mel_filter_coefs[38][16] = 16'h0000;
	mel_filter_coefs[38][17] = 16'h0000;
	mel_filter_coefs[38][18] = 16'h0000;
	mel_filter_coefs[38][19] = 16'h0000;
	mel_filter_coefs[38][20] = 16'h0000;
	mel_filter_coefs[38][21] = 16'h0000;
	mel_filter_coefs[38][22] = 16'h0000;
	mel_filter_coefs[38][23] = 16'h0000;
	mel_filter_coefs[38][24] = 16'h0000;
	mel_filter_coefs[38][25] = 16'h0000;
	mel_filter_coefs[38][26] = 16'h0000;
	mel_filter_coefs[38][27] = 16'h0000;
	mel_filter_coefs[38][28] = 16'h0000;
	mel_filter_coefs[38][29] = 16'h0000;
	mel_filter_coefs[38][30] = 16'h0000;
	mel_filter_coefs[38][31] = 16'h0000;
	mel_filter_coefs[38][32] = 16'h0000;
	mel_filter_coefs[38][33] = 16'h0000;
	mel_filter_coefs[38][34] = 16'h0000;
	mel_filter_coefs[38][35] = 16'h0000;
	mel_filter_coefs[38][36] = 16'h0000;
	mel_filter_coefs[38][37] = 16'h0000;
	mel_filter_coefs[38][38] = 16'h0000;
	mel_filter_coefs[38][39] = 16'h0000;
	mel_filter_coefs[38][40] = 16'h0000;
	mel_filter_coefs[38][41] = 16'h0000;
	mel_filter_coefs[38][42] = 16'h0000;
	mel_filter_coefs[38][43] = 16'h0000;
	mel_filter_coefs[38][44] = 16'h0000;
	mel_filter_coefs[38][45] = 16'h0000;
	mel_filter_coefs[38][46] = 16'h0000;
	mel_filter_coefs[38][47] = 16'h0000;
	mel_filter_coefs[38][48] = 16'h0000;
	mel_filter_coefs[38][49] = 16'h0000;
	mel_filter_coefs[38][50] = 16'h0000;
	mel_filter_coefs[38][51] = 16'h0000;
	mel_filter_coefs[38][52] = 16'h0000;
	mel_filter_coefs[38][53] = 16'h0000;
	mel_filter_coefs[38][54] = 16'h0000;
	mel_filter_coefs[38][55] = 16'h0000;
	mel_filter_coefs[38][56] = 16'h0000;
	mel_filter_coefs[38][57] = 16'h0000;
	mel_filter_coefs[38][58] = 16'h0000;
	mel_filter_coefs[38][59] = 16'h0000;
	mel_filter_coefs[38][60] = 16'h0000;
	mel_filter_coefs[38][61] = 16'h0000;
	mel_filter_coefs[38][62] = 16'h0000;
	mel_filter_coefs[38][63] = 16'h0000;
	mel_filter_coefs[38][64] = 16'h0000;
	mel_filter_coefs[38][65] = 16'h0000;
	mel_filter_coefs[38][66] = 16'h0000;
	mel_filter_coefs[38][67] = 16'h0000;
	mel_filter_coefs[38][68] = 16'h0000;
	mel_filter_coefs[38][69] = 16'h0000;
	mel_filter_coefs[38][70] = 16'h0000;
	mel_filter_coefs[38][71] = 16'h0000;
	mel_filter_coefs[38][72] = 16'h0000;
	mel_filter_coefs[38][73] = 16'h0000;
	mel_filter_coefs[38][74] = 16'h0000;
	mel_filter_coefs[38][75] = 16'h0000;
	mel_filter_coefs[38][76] = 16'h0000;
	mel_filter_coefs[38][77] = 16'h0000;
	mel_filter_coefs[38][78] = 16'h0000;
	mel_filter_coefs[38][79] = 16'h0000;
	mel_filter_coefs[38][80] = 16'h0000;
	mel_filter_coefs[38][81] = 16'h0000;
	mel_filter_coefs[38][82] = 16'h0000;
	mel_filter_coefs[38][83] = 16'h0000;
	mel_filter_coefs[38][84] = 16'h0000;
	mel_filter_coefs[38][85] = 16'h0000;
	mel_filter_coefs[38][86] = 16'h0000;
	mel_filter_coefs[38][87] = 16'h0000;
	mel_filter_coefs[38][88] = 16'h0000;
	mel_filter_coefs[38][89] = 16'h0000;
	mel_filter_coefs[38][90] = 16'h0000;
	mel_filter_coefs[38][91] = 16'h0000;
	mel_filter_coefs[38][92] = 16'h0000;
	mel_filter_coefs[38][93] = 16'h0000;
	mel_filter_coefs[38][94] = 16'h0000;
	mel_filter_coefs[38][95] = 16'h0000;
	mel_filter_coefs[38][96] = 16'h0000;
	mel_filter_coefs[38][97] = 16'h0000;
	mel_filter_coefs[38][98] = 16'h0000;
	mel_filter_coefs[38][99] = 16'h0000;
	mel_filter_coefs[38][100] = 16'h0000;
	mel_filter_coefs[38][101] = 16'h0000;
	mel_filter_coefs[38][102] = 16'h0000;
	mel_filter_coefs[38][103] = 16'h0000;
	mel_filter_coefs[38][104] = 16'h0000;
	mel_filter_coefs[38][105] = 16'h0000;
	mel_filter_coefs[38][106] = 16'h0000;
	mel_filter_coefs[38][107] = 16'h0000;
	mel_filter_coefs[38][108] = 16'h0000;
	mel_filter_coefs[38][109] = 16'h0000;
	mel_filter_coefs[38][110] = 16'h0000;
	mel_filter_coefs[38][111] = 16'h0000;
	mel_filter_coefs[38][112] = 16'h0000;
	mel_filter_coefs[38][113] = 16'h0000;
	mel_filter_coefs[38][114] = 16'h0000;
	mel_filter_coefs[38][115] = 16'h0000;
	mel_filter_coefs[38][116] = 16'h0000;
	mel_filter_coefs[38][117] = 16'h0000;
	mel_filter_coefs[38][118] = 16'h0000;
	mel_filter_coefs[38][119] = 16'h0000;
	mel_filter_coefs[38][120] = 16'h0000;
	mel_filter_coefs[38][121] = 16'h0000;
	mel_filter_coefs[38][122] = 16'h0000;
	mel_filter_coefs[38][123] = 16'h0000;
	mel_filter_coefs[38][124] = 16'h0000;
	mel_filter_coefs[38][125] = 16'h0000;
	mel_filter_coefs[38][126] = 16'h0000;
	mel_filter_coefs[38][127] = 16'h0000;
	mel_filter_coefs[38][128] = 16'h0000;
	mel_filter_coefs[38][129] = 16'h0000;
	mel_filter_coefs[38][130] = 16'h0000;
	mel_filter_coefs[38][131] = 16'h0000;
	mel_filter_coefs[38][132] = 16'h0000;
	mel_filter_coefs[38][133] = 16'h0000;
	mel_filter_coefs[38][134] = 16'h0000;
	mel_filter_coefs[38][135] = 16'h0000;
	mel_filter_coefs[38][136] = 16'h0000;
	mel_filter_coefs[38][137] = 16'h0000;
	mel_filter_coefs[38][138] = 16'h0000;
	mel_filter_coefs[38][139] = 16'h0000;
	mel_filter_coefs[38][140] = 16'h0000;
	mel_filter_coefs[38][141] = 16'h0000;
	mel_filter_coefs[38][142] = 16'h0000;
	mel_filter_coefs[38][143] = 16'h0000;
	mel_filter_coefs[38][144] = 16'h0000;
	mel_filter_coefs[38][145] = 16'h0000;
	mel_filter_coefs[38][146] = 16'h0000;
	mel_filter_coefs[38][147] = 16'h0000;
	mel_filter_coefs[38][148] = 16'h0000;
	mel_filter_coefs[38][149] = 16'h0000;
	mel_filter_coefs[38][150] = 16'h0000;
	mel_filter_coefs[38][151] = 16'h0000;
	mel_filter_coefs[38][152] = 16'h0000;
	mel_filter_coefs[38][153] = 16'h0000;
	mel_filter_coefs[38][154] = 16'h0000;
	mel_filter_coefs[38][155] = 16'h0000;
	mel_filter_coefs[38][156] = 16'h0000;
	mel_filter_coefs[38][157] = 16'h0000;
	mel_filter_coefs[38][158] = 16'h0000;
	mel_filter_coefs[38][159] = 16'h0000;
	mel_filter_coefs[38][160] = 16'h0000;
	mel_filter_coefs[38][161] = 16'h0000;
	mel_filter_coefs[38][162] = 16'h0000;
	mel_filter_coefs[38][163] = 16'h0000;
	mel_filter_coefs[38][164] = 16'h0000;
	mel_filter_coefs[38][165] = 16'h0000;
	mel_filter_coefs[38][166] = 16'h0000;
	mel_filter_coefs[38][167] = 16'h0000;
	mel_filter_coefs[38][168] = 16'h0000;
	mel_filter_coefs[38][169] = 16'h0000;
	mel_filter_coefs[38][170] = 16'h0000;
	mel_filter_coefs[38][171] = 16'h0000;
	mel_filter_coefs[38][172] = 16'h0000;
	mel_filter_coefs[38][173] = 16'h0000;
	mel_filter_coefs[38][174] = 16'h0000;
	mel_filter_coefs[38][175] = 16'h0000;
	mel_filter_coefs[38][176] = 16'h0000;
	mel_filter_coefs[38][177] = 16'h0000;
	mel_filter_coefs[38][178] = 16'h0000;
	mel_filter_coefs[38][179] = 16'h0000;
	mel_filter_coefs[38][180] = 16'h0000;
	mel_filter_coefs[38][181] = 16'h0000;
	mel_filter_coefs[38][182] = 16'h0000;
	mel_filter_coefs[38][183] = 16'h0000;
	mel_filter_coefs[38][184] = 16'h0000;
	mel_filter_coefs[38][185] = 16'h0000;
	mel_filter_coefs[38][186] = 16'h0000;
	mel_filter_coefs[38][187] = 16'h0000;
	mel_filter_coefs[38][188] = 16'h0000;
	mel_filter_coefs[38][189] = 16'h0000;
	mel_filter_coefs[38][190] = 16'h0000;
	mel_filter_coefs[38][191] = 16'h0000;
	mel_filter_coefs[38][192] = 16'h0000;
	mel_filter_coefs[38][193] = 16'h0000;
	mel_filter_coefs[38][194] = 16'h0000;
	mel_filter_coefs[38][195] = 16'h0000;
	mel_filter_coefs[38][196] = 16'h0000;
	mel_filter_coefs[38][197] = 16'h0000;
	mel_filter_coefs[38][198] = 16'h0000;
	mel_filter_coefs[38][199] = 16'h0000;
	mel_filter_coefs[38][200] = 16'h0000;
	mel_filter_coefs[38][201] = 16'h0000;
	mel_filter_coefs[38][202] = 16'h0000;
	mel_filter_coefs[38][203] = 16'h0000;
	mel_filter_coefs[38][204] = 16'h0000;
	mel_filter_coefs[38][205] = 16'h0000;
	mel_filter_coefs[38][206] = 16'h0000;
	mel_filter_coefs[38][207] = 16'h0000;
	mel_filter_coefs[38][208] = 16'h0000;
	mel_filter_coefs[38][209] = 16'h0619;
	mel_filter_coefs[38][210] = 16'h0EDA;
	mel_filter_coefs[38][211] = 16'h179C;
	mel_filter_coefs[38][212] = 16'h205D;
	mel_filter_coefs[38][213] = 16'h291E;
	mel_filter_coefs[38][214] = 16'h31E0;
	mel_filter_coefs[38][215] = 16'h3AA1;
	mel_filter_coefs[38][216] = 16'h4363;
	mel_filter_coefs[38][217] = 16'h4C24;
	mel_filter_coefs[38][218] = 16'h54E6;
	mel_filter_coefs[38][219] = 16'h5DA7;
	mel_filter_coefs[38][220] = 16'h6669;
	mel_filter_coefs[38][221] = 16'h6F2A;
	mel_filter_coefs[38][222] = 16'h77EC;
	mel_filter_coefs[38][223] = 16'h7F5D;
	mel_filter_coefs[38][224] = 16'h7722;
	mel_filter_coefs[38][225] = 16'h6EE6;
	mel_filter_coefs[38][226] = 16'h66AA;
	mel_filter_coefs[38][227] = 16'h5E6E;
	mel_filter_coefs[38][228] = 16'h5632;
	mel_filter_coefs[38][229] = 16'h4DF6;
	mel_filter_coefs[38][230] = 16'h45BB;
	mel_filter_coefs[38][231] = 16'h3D7F;
	mel_filter_coefs[38][232] = 16'h3543;
	mel_filter_coefs[38][233] = 16'h2D07;
	mel_filter_coefs[38][234] = 16'h24CB;
	mel_filter_coefs[38][235] = 16'h1C8F;
	mel_filter_coefs[38][236] = 16'h1454;
	mel_filter_coefs[38][237] = 16'h0C18;
	mel_filter_coefs[38][238] = 16'h03DC;
	mel_filter_coefs[38][239] = 16'h0000;
	mel_filter_coefs[38][240] = 16'h0000;
	mel_filter_coefs[38][241] = 16'h0000;
	mel_filter_coefs[38][242] = 16'h0000;
	mel_filter_coefs[38][243] = 16'h0000;
	mel_filter_coefs[38][244] = 16'h0000;
	mel_filter_coefs[38][245] = 16'h0000;
	mel_filter_coefs[38][246] = 16'h0000;
	mel_filter_coefs[38][247] = 16'h0000;
	mel_filter_coefs[38][248] = 16'h0000;
	mel_filter_coefs[38][249] = 16'h0000;
	mel_filter_coefs[38][250] = 16'h0000;
	mel_filter_coefs[38][251] = 16'h0000;
	mel_filter_coefs[38][252] = 16'h0000;
	mel_filter_coefs[38][253] = 16'h0000;
	mel_filter_coefs[38][254] = 16'h0000;
	mel_filter_coefs[38][255] = 16'h0000;
	mel_filter_coefs[39][0] = 16'h0000;
	mel_filter_coefs[39][1] = 16'h0000;
	mel_filter_coefs[39][2] = 16'h0000;
	mel_filter_coefs[39][3] = 16'h0000;
	mel_filter_coefs[39][4] = 16'h0000;
	mel_filter_coefs[39][5] = 16'h0000;
	mel_filter_coefs[39][6] = 16'h0000;
	mel_filter_coefs[39][7] = 16'h0000;
	mel_filter_coefs[39][8] = 16'h0000;
	mel_filter_coefs[39][9] = 16'h0000;
	mel_filter_coefs[39][10] = 16'h0000;
	mel_filter_coefs[39][11] = 16'h0000;
	mel_filter_coefs[39][12] = 16'h0000;
	mel_filter_coefs[39][13] = 16'h0000;
	mel_filter_coefs[39][14] = 16'h0000;
	mel_filter_coefs[39][15] = 16'h0000;
	mel_filter_coefs[39][16] = 16'h0000;
	mel_filter_coefs[39][17] = 16'h0000;
	mel_filter_coefs[39][18] = 16'h0000;
	mel_filter_coefs[39][19] = 16'h0000;
	mel_filter_coefs[39][20] = 16'h0000;
	mel_filter_coefs[39][21] = 16'h0000;
	mel_filter_coefs[39][22] = 16'h0000;
	mel_filter_coefs[39][23] = 16'h0000;
	mel_filter_coefs[39][24] = 16'h0000;
	mel_filter_coefs[39][25] = 16'h0000;
	mel_filter_coefs[39][26] = 16'h0000;
	mel_filter_coefs[39][27] = 16'h0000;
	mel_filter_coefs[39][28] = 16'h0000;
	mel_filter_coefs[39][29] = 16'h0000;
	mel_filter_coefs[39][30] = 16'h0000;
	mel_filter_coefs[39][31] = 16'h0000;
	mel_filter_coefs[39][32] = 16'h0000;
	mel_filter_coefs[39][33] = 16'h0000;
	mel_filter_coefs[39][34] = 16'h0000;
	mel_filter_coefs[39][35] = 16'h0000;
	mel_filter_coefs[39][36] = 16'h0000;
	mel_filter_coefs[39][37] = 16'h0000;
	mel_filter_coefs[39][38] = 16'h0000;
	mel_filter_coefs[39][39] = 16'h0000;
	mel_filter_coefs[39][40] = 16'h0000;
	mel_filter_coefs[39][41] = 16'h0000;
	mel_filter_coefs[39][42] = 16'h0000;
	mel_filter_coefs[39][43] = 16'h0000;
	mel_filter_coefs[39][44] = 16'h0000;
	mel_filter_coefs[39][45] = 16'h0000;
	mel_filter_coefs[39][46] = 16'h0000;
	mel_filter_coefs[39][47] = 16'h0000;
	mel_filter_coefs[39][48] = 16'h0000;
	mel_filter_coefs[39][49] = 16'h0000;
	mel_filter_coefs[39][50] = 16'h0000;
	mel_filter_coefs[39][51] = 16'h0000;
	mel_filter_coefs[39][52] = 16'h0000;
	mel_filter_coefs[39][53] = 16'h0000;
	mel_filter_coefs[39][54] = 16'h0000;
	mel_filter_coefs[39][55] = 16'h0000;
	mel_filter_coefs[39][56] = 16'h0000;
	mel_filter_coefs[39][57] = 16'h0000;
	mel_filter_coefs[39][58] = 16'h0000;
	mel_filter_coefs[39][59] = 16'h0000;
	mel_filter_coefs[39][60] = 16'h0000;
	mel_filter_coefs[39][61] = 16'h0000;
	mel_filter_coefs[39][62] = 16'h0000;
	mel_filter_coefs[39][63] = 16'h0000;
	mel_filter_coefs[39][64] = 16'h0000;
	mel_filter_coefs[39][65] = 16'h0000;
	mel_filter_coefs[39][66] = 16'h0000;
	mel_filter_coefs[39][67] = 16'h0000;
	mel_filter_coefs[39][68] = 16'h0000;
	mel_filter_coefs[39][69] = 16'h0000;
	mel_filter_coefs[39][70] = 16'h0000;
	mel_filter_coefs[39][71] = 16'h0000;
	mel_filter_coefs[39][72] = 16'h0000;
	mel_filter_coefs[39][73] = 16'h0000;
	mel_filter_coefs[39][74] = 16'h0000;
	mel_filter_coefs[39][75] = 16'h0000;
	mel_filter_coefs[39][76] = 16'h0000;
	mel_filter_coefs[39][77] = 16'h0000;
	mel_filter_coefs[39][78] = 16'h0000;
	mel_filter_coefs[39][79] = 16'h0000;
	mel_filter_coefs[39][80] = 16'h0000;
	mel_filter_coefs[39][81] = 16'h0000;
	mel_filter_coefs[39][82] = 16'h0000;
	mel_filter_coefs[39][83] = 16'h0000;
	mel_filter_coefs[39][84] = 16'h0000;
	mel_filter_coefs[39][85] = 16'h0000;
	mel_filter_coefs[39][86] = 16'h0000;
	mel_filter_coefs[39][87] = 16'h0000;
	mel_filter_coefs[39][88] = 16'h0000;
	mel_filter_coefs[39][89] = 16'h0000;
	mel_filter_coefs[39][90] = 16'h0000;
	mel_filter_coefs[39][91] = 16'h0000;
	mel_filter_coefs[39][92] = 16'h0000;
	mel_filter_coefs[39][93] = 16'h0000;
	mel_filter_coefs[39][94] = 16'h0000;
	mel_filter_coefs[39][95] = 16'h0000;
	mel_filter_coefs[39][96] = 16'h0000;
	mel_filter_coefs[39][97] = 16'h0000;
	mel_filter_coefs[39][98] = 16'h0000;
	mel_filter_coefs[39][99] = 16'h0000;
	mel_filter_coefs[39][100] = 16'h0000;
	mel_filter_coefs[39][101] = 16'h0000;
	mel_filter_coefs[39][102] = 16'h0000;
	mel_filter_coefs[39][103] = 16'h0000;
	mel_filter_coefs[39][104] = 16'h0000;
	mel_filter_coefs[39][105] = 16'h0000;
	mel_filter_coefs[39][106] = 16'h0000;
	mel_filter_coefs[39][107] = 16'h0000;
	mel_filter_coefs[39][108] = 16'h0000;
	mel_filter_coefs[39][109] = 16'h0000;
	mel_filter_coefs[39][110] = 16'h0000;
	mel_filter_coefs[39][111] = 16'h0000;
	mel_filter_coefs[39][112] = 16'h0000;
	mel_filter_coefs[39][113] = 16'h0000;
	mel_filter_coefs[39][114] = 16'h0000;
	mel_filter_coefs[39][115] = 16'h0000;
	mel_filter_coefs[39][116] = 16'h0000;
	mel_filter_coefs[39][117] = 16'h0000;
	mel_filter_coefs[39][118] = 16'h0000;
	mel_filter_coefs[39][119] = 16'h0000;
	mel_filter_coefs[39][120] = 16'h0000;
	mel_filter_coefs[39][121] = 16'h0000;
	mel_filter_coefs[39][122] = 16'h0000;
	mel_filter_coefs[39][123] = 16'h0000;
	mel_filter_coefs[39][124] = 16'h0000;
	mel_filter_coefs[39][125] = 16'h0000;
	mel_filter_coefs[39][126] = 16'h0000;
	mel_filter_coefs[39][127] = 16'h0000;
	mel_filter_coefs[39][128] = 16'h0000;
	mel_filter_coefs[39][129] = 16'h0000;
	mel_filter_coefs[39][130] = 16'h0000;
	mel_filter_coefs[39][131] = 16'h0000;
	mel_filter_coefs[39][132] = 16'h0000;
	mel_filter_coefs[39][133] = 16'h0000;
	mel_filter_coefs[39][134] = 16'h0000;
	mel_filter_coefs[39][135] = 16'h0000;
	mel_filter_coefs[39][136] = 16'h0000;
	mel_filter_coefs[39][137] = 16'h0000;
	mel_filter_coefs[39][138] = 16'h0000;
	mel_filter_coefs[39][139] = 16'h0000;
	mel_filter_coefs[39][140] = 16'h0000;
	mel_filter_coefs[39][141] = 16'h0000;
	mel_filter_coefs[39][142] = 16'h0000;
	mel_filter_coefs[39][143] = 16'h0000;
	mel_filter_coefs[39][144] = 16'h0000;
	mel_filter_coefs[39][145] = 16'h0000;
	mel_filter_coefs[39][146] = 16'h0000;
	mel_filter_coefs[39][147] = 16'h0000;
	mel_filter_coefs[39][148] = 16'h0000;
	mel_filter_coefs[39][149] = 16'h0000;
	mel_filter_coefs[39][150] = 16'h0000;
	mel_filter_coefs[39][151] = 16'h0000;
	mel_filter_coefs[39][152] = 16'h0000;
	mel_filter_coefs[39][153] = 16'h0000;
	mel_filter_coefs[39][154] = 16'h0000;
	mel_filter_coefs[39][155] = 16'h0000;
	mel_filter_coefs[39][156] = 16'h0000;
	mel_filter_coefs[39][157] = 16'h0000;
	mel_filter_coefs[39][158] = 16'h0000;
	mel_filter_coefs[39][159] = 16'h0000;
	mel_filter_coefs[39][160] = 16'h0000;
	mel_filter_coefs[39][161] = 16'h0000;
	mel_filter_coefs[39][162] = 16'h0000;
	mel_filter_coefs[39][163] = 16'h0000;
	mel_filter_coefs[39][164] = 16'h0000;
	mel_filter_coefs[39][165] = 16'h0000;
	mel_filter_coefs[39][166] = 16'h0000;
	mel_filter_coefs[39][167] = 16'h0000;
	mel_filter_coefs[39][168] = 16'h0000;
	mel_filter_coefs[39][169] = 16'h0000;
	mel_filter_coefs[39][170] = 16'h0000;
	mel_filter_coefs[39][171] = 16'h0000;
	mel_filter_coefs[39][172] = 16'h0000;
	mel_filter_coefs[39][173] = 16'h0000;
	mel_filter_coefs[39][174] = 16'h0000;
	mel_filter_coefs[39][175] = 16'h0000;
	mel_filter_coefs[39][176] = 16'h0000;
	mel_filter_coefs[39][177] = 16'h0000;
	mel_filter_coefs[39][178] = 16'h0000;
	mel_filter_coefs[39][179] = 16'h0000;
	mel_filter_coefs[39][180] = 16'h0000;
	mel_filter_coefs[39][181] = 16'h0000;
	mel_filter_coefs[39][182] = 16'h0000;
	mel_filter_coefs[39][183] = 16'h0000;
	mel_filter_coefs[39][184] = 16'h0000;
	mel_filter_coefs[39][185] = 16'h0000;
	mel_filter_coefs[39][186] = 16'h0000;
	mel_filter_coefs[39][187] = 16'h0000;
	mel_filter_coefs[39][188] = 16'h0000;
	mel_filter_coefs[39][189] = 16'h0000;
	mel_filter_coefs[39][190] = 16'h0000;
	mel_filter_coefs[39][191] = 16'h0000;
	mel_filter_coefs[39][192] = 16'h0000;
	mel_filter_coefs[39][193] = 16'h0000;
	mel_filter_coefs[39][194] = 16'h0000;
	mel_filter_coefs[39][195] = 16'h0000;
	mel_filter_coefs[39][196] = 16'h0000;
	mel_filter_coefs[39][197] = 16'h0000;
	mel_filter_coefs[39][198] = 16'h0000;
	mel_filter_coefs[39][199] = 16'h0000;
	mel_filter_coefs[39][200] = 16'h0000;
	mel_filter_coefs[39][201] = 16'h0000;
	mel_filter_coefs[39][202] = 16'h0000;
	mel_filter_coefs[39][203] = 16'h0000;
	mel_filter_coefs[39][204] = 16'h0000;
	mel_filter_coefs[39][205] = 16'h0000;
	mel_filter_coefs[39][206] = 16'h0000;
	mel_filter_coefs[39][207] = 16'h0000;
	mel_filter_coefs[39][208] = 16'h0000;
	mel_filter_coefs[39][209] = 16'h0000;
	mel_filter_coefs[39][210] = 16'h0000;
	mel_filter_coefs[39][211] = 16'h0000;
	mel_filter_coefs[39][212] = 16'h0000;
	mel_filter_coefs[39][213] = 16'h0000;
	mel_filter_coefs[39][214] = 16'h0000;
	mel_filter_coefs[39][215] = 16'h0000;
	mel_filter_coefs[39][216] = 16'h0000;
	mel_filter_coefs[39][217] = 16'h0000;
	mel_filter_coefs[39][218] = 16'h0000;
	mel_filter_coefs[39][219] = 16'h0000;
	mel_filter_coefs[39][220] = 16'h0000;
	mel_filter_coefs[39][221] = 16'h0000;
	mel_filter_coefs[39][222] = 16'h0000;
	mel_filter_coefs[39][223] = 16'h00A3;
	mel_filter_coefs[39][224] = 16'h08DE;
	mel_filter_coefs[39][225] = 16'h111A;
	mel_filter_coefs[39][226] = 16'h1956;
	mel_filter_coefs[39][227] = 16'h2192;
	mel_filter_coefs[39][228] = 16'h29CE;
	mel_filter_coefs[39][229] = 16'h320A;
	mel_filter_coefs[39][230] = 16'h3A45;
	mel_filter_coefs[39][231] = 16'h4281;
	mel_filter_coefs[39][232] = 16'h4ABD;
	mel_filter_coefs[39][233] = 16'h52F9;
	mel_filter_coefs[39][234] = 16'h5B35;
	mel_filter_coefs[39][235] = 16'h6371;
	mel_filter_coefs[39][236] = 16'h6BAC;
	mel_filter_coefs[39][237] = 16'h73E8;
	mel_filter_coefs[39][238] = 16'h7C24;
	mel_filter_coefs[39][239] = 16'h7BE3;
	mel_filter_coefs[39][240] = 16'h7425;
	mel_filter_coefs[39][241] = 16'h6C66;
	mel_filter_coefs[39][242] = 16'h64A8;
	mel_filter_coefs[39][243] = 16'h5CEA;
	mel_filter_coefs[39][244] = 16'h552C;
	mel_filter_coefs[39][245] = 16'h4D6E;
	mel_filter_coefs[39][246] = 16'h45B0;
	mel_filter_coefs[39][247] = 16'h3DF1;
	mel_filter_coefs[39][248] = 16'h3633;
	mel_filter_coefs[39][249] = 16'h2E75;
	mel_filter_coefs[39][250] = 16'h26B7;
	mel_filter_coefs[39][251] = 16'h1EF9;
	mel_filter_coefs[39][252] = 16'h173B;
	mel_filter_coefs[39][253] = 16'h0F7C;
	mel_filter_coefs[39][254] = 16'h07BE;
	mel_filter_coefs[39][255] = 16'h0000;

	end

    // Mel-scale filterbank computation
    integer i;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            mel_filter_cnt <= 0;
            dft_point_cnt <= 0;
            mel_fbank_out <= 0;
            mel_fbank_valid <= 0;
            for (i = 0; i < NUM_MEL_FILTERS; i = i + 1) begin
                mel_accumulators[i] <= 0;
            end
        end else begin
            if (dft_valid) begin
                // Multiply DFT output with the corresponding filter coefficient
                mel_accumulators[mel_filter_cnt] <= mel_accumulators[mel_filter_cnt] +
                    (dft_out * mel_filter_coefs[mel_filter_cnt][dft_point_cnt]);

                // Increment DFT point counter
                if (dft_point_cnt == NUM_DFT_POINTS - 1) begin
                    dft_point_cnt <= 0;

                    // Increment mel-scale filter counter
                    if (mel_filter_cnt == NUM_MEL_FILTERS - 1) begin
                        mel_filter_cnt <= 0;

                        // Output the accumulated filterbank energies
                        mel_fbank_out <= mel_accumulators[NUM_MEL_FILTERS - 1];
                        mel_fbank_valid <= 1;

                        // Reset the accumulators for the next frame
                        for (i = 0; i < NUM_MEL_FILTERS; i = i + 1) begin
                            mel_accumulators[i] <= 0;
                        end
                    end else begin
                        mel_filter_cnt <= mel_filter_cnt + 1;
                        mel_fbank_out <= 0;
                        mel_fbank_valid <= 0;
                    end
                end else begin
                    dft_point_cnt <= dft_point_cnt + 1;
                    mel_fbank_out <= 0;
                    mel_fbank_valid <= 0;
                end
            end else begin
                mel_fbank_out <= 0;
                mel_fbank_valid <= 0;
            end
        end
    end

endmodule

`endif
